magic
tech sky130A
timestamp 1645554640
<< error_p >>
rect 900 1488 1338 1498
rect 1381 1488 1499 1498
rect 900 912 912 1488
rect 900 900 1338 912
rect 1381 900 1499 912
<< metal4 >>
rect -600 1498 1500 1500
rect -600 900 900 1498
rect 1338 1380 1381 1498
rect 1499 1380 1500 1498
rect 1338 1338 1500 1380
rect 1338 1220 1381 1338
rect 1499 1220 1500 1338
rect 1338 1178 1500 1220
rect 1338 1060 1381 1178
rect 1499 1060 1500 1178
rect 1338 1018 1500 1060
rect 1338 900 1381 1018
rect 1499 900 1500 1018
<< via4 >>
rect 900 900 1338 1498
rect 1381 1380 1499 1498
rect 1381 1220 1499 1338
rect 1381 1060 1499 1178
rect 1381 900 1499 1018
<< metal5 >>
rect 0 14400 15000 15000
rect 0 13500 14100 14100
rect 0 600 600 13500
rect 13500 1500 14100 13500
rect 900 1498 14100 1500
rect 1338 1380 1381 1498
rect 1499 1380 14100 1498
rect 1338 1338 14100 1380
rect 1338 1220 1381 1338
rect 1499 1220 14100 1338
rect 1338 1178 14100 1220
rect 1338 1060 1381 1178
rect 1499 1060 14100 1178
rect 1338 1018 14100 1060
rect 1338 900 1381 1018
rect 1499 900 14100 1018
rect 14400 600 15000 14400
rect 0 0 15000 600
<< end >>
