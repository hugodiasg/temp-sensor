magic
tech sky130A
magscale 1 2
timestamp 1643668240
<< metal3 >>
rect -2125 2047 2124 2075
rect -2125 -2047 2040 2047
rect 2104 -2047 2124 2047
rect -2125 -2075 2124 -2047
<< via3 >>
rect 2040 -2047 2104 2047
<< mimcap >>
rect -2025 1935 1925 1975
rect -2025 -1935 -1985 1935
rect 1885 -1935 1925 1935
rect -2025 -1975 1925 -1935
<< mimcapcontact >>
rect -1985 -1935 1885 1935
<< metal4 >>
rect 2024 2047 2120 2063
rect -1986 1935 1886 1936
rect -1986 -1935 -1985 1935
rect 1885 -1935 1886 1935
rect -1986 -1936 1886 -1935
rect 2024 -2047 2040 2047
rect 2104 -2047 2120 2047
rect 2024 -2063 2120 -2047
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -2125 -2075 2025 2075
string parameters w 19.75 l 19.75 val 795.135 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
