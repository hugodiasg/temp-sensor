magic
tech sky130A
magscale 1 2
timestamp 1656776172
<< nwell >>
rect -1560 -4780 -168 -3942
<< pmos >>
rect -1364 -4561 -364 -4161
<< pdiff >>
rect -1422 -4173 -1364 -4161
rect -1422 -4549 -1410 -4173
rect -1376 -4549 -1364 -4173
rect -1422 -4561 -1364 -4549
rect -364 -4173 -306 -4161
rect -364 -4549 -352 -4173
rect -318 -4549 -306 -4173
rect -364 -4561 -306 -4549
<< pdiffc >>
rect -1410 -4549 -1376 -4173
rect -352 -4549 -318 -4173
<< psubdiff >>
rect 2820 -4860 2920 -4836
rect 2820 -4984 2920 -4960
<< nsubdiff >>
rect -1524 -4012 -1428 -3978
rect -300 -4012 -204 -3978
rect -1524 -4074 -1490 -4012
rect -238 -4074 -204 -4012
rect -1524 -4710 -1490 -4648
rect -238 -4710 -204 -4648
rect -1524 -4744 -1428 -4710
rect -300 -4744 -204 -4710
<< psubdiffcont >>
rect 2820 -4960 2920 -4860
<< nsubdiffcont >>
rect -1428 -4012 -300 -3978
rect -1524 -4648 -1490 -4074
rect -238 -4648 -204 -4074
rect -1428 -4744 -300 -4710
<< poly >>
rect -1364 -4080 -364 -4064
rect -1364 -4114 -1348 -4080
rect -380 -4114 -364 -4080
rect -1364 -4161 -364 -4114
rect -1364 -4608 -364 -4561
rect -1364 -4642 -1348 -4608
rect -380 -4642 -364 -4608
rect -1364 -4658 -364 -4642
<< polycont >>
rect -1348 -4114 -380 -4080
rect -1348 -4642 -380 -4608
<< locali >>
rect -1524 -4012 -1428 -3978
rect -300 -4012 -204 -3978
rect -1524 -4074 -1490 -4012
rect -238 -4074 -204 -4012
rect -1364 -4114 -1348 -4080
rect -380 -4114 -364 -4080
rect -1410 -4173 -1376 -4157
rect -1410 -4565 -1376 -4549
rect -352 -4173 -318 -4157
rect -352 -4565 -318 -4549
rect -1364 -4642 -1348 -4608
rect -380 -4642 -364 -4608
rect -1524 -4710 -1490 -4648
rect -238 -4710 -204 -4648
rect -1524 -4744 -1428 -4710
rect -300 -4744 -204 -4710
<< viali >>
rect 2820 -4860 2920 -4840
rect 2820 -4960 2920 -4860
rect 2820 -4980 2920 -4960
<< metal1 >>
rect -1840 -1380 -1640 -940
rect -240 -1200 -40 -940
rect -2100 -1560 -1400 -1380
rect -1580 -2240 -1400 -1560
rect -240 -1400 980 -1200
rect 1840 -1380 3200 -1300
rect -240 -1840 -40 -1400
rect 800 -1480 980 -1400
rect 1180 -1440 1760 -1380
rect 800 -1660 1180 -1480
rect 1380 -1580 1760 -1440
rect 1840 -1440 1860 -1380
rect 1920 -1420 2460 -1380
rect 1920 -1440 1940 -1420
rect 1840 -1460 1940 -1440
rect 1400 -1600 1760 -1580
rect 104 -1840 296 -1838
rect -360 -1850 296 -1840
rect -367 -1901 296 -1850
rect -360 -2220 280 -1901
rect 480 -2160 580 -2140
rect 480 -2220 500 -2160
rect 560 -2220 580 -2160
rect 480 -2240 580 -2220
rect -1000 -2300 -740 -2280
rect 360 -2300 420 -2280
rect -2360 -4780 -2140 -4500
rect -1280 -4780 -440 -2300
rect 320 -2540 460 -2300
rect -140 -2660 460 -2540
rect 1200 -2640 1360 -2320
rect -140 -4780 40 -2660
rect 500 -2700 1360 -2640
rect 300 -2760 1360 -2700
rect 300 -2940 500 -2760
rect 220 -3000 320 -2980
rect 1340 -3000 1440 -2980
rect 120 -3060 240 -3000
rect 300 -3060 320 -3000
rect 220 -3080 320 -3060
rect 520 -3700 1140 -3000
rect 1340 -3060 1360 -3000
rect 1420 -3060 1440 -3000
rect 1340 -3080 1440 -3060
rect 520 -3760 1160 -3700
rect 520 -4580 1140 -3760
rect 1640 -4580 1760 -1600
rect 1840 -1820 1940 -1800
rect 1840 -1880 1860 -1820
rect 1920 -1880 1940 -1820
rect 1840 -1900 1940 -1880
rect 1840 -2240 1940 -2200
rect 1840 -2300 1860 -2240
rect 1920 -2300 1940 -2240
rect 1840 -2660 1940 -2640
rect 1840 -2720 1860 -2660
rect 1920 -2720 1940 -2660
rect 1840 -2740 1940 -2720
rect 1840 -3060 1940 -3040
rect 1840 -3120 1860 -3060
rect 1920 -3120 1940 -3060
rect 1840 -3140 1940 -3120
rect 1840 -3500 1940 -3480
rect 1840 -3560 1860 -3500
rect 1920 -3560 1940 -3500
rect 1840 -3580 1940 -3560
rect 1840 -3900 1940 -3880
rect 1840 -3960 1860 -3900
rect 1920 -3960 1940 -3900
rect 1840 -3980 1940 -3960
rect 1840 -4320 1940 -4300
rect 1840 -4380 1860 -4320
rect 1920 -4380 1940 -4320
rect 1840 -4400 1940 -4380
rect 1180 -4720 1240 -4620
rect 1320 -4720 1380 -4620
rect 1180 -4780 1380 -4720
rect -2360 -4920 1380 -4780
rect 2020 -4800 2140 -1460
rect 2240 -4600 2360 -1420
rect 2440 -1440 2460 -1420
rect 2520 -1420 3060 -1380
rect 2520 -1440 2540 -1420
rect 2440 -1460 2540 -1440
rect 3040 -1440 3060 -1420
rect 3120 -1420 3200 -1380
rect 3120 -1440 3142 -1420
rect 3040 -1460 3142 -1440
rect 2440 -1820 2540 -1780
rect 2440 -1880 2460 -1820
rect 2520 -1880 2540 -1820
rect 2440 -1900 2540 -1880
rect 2440 -2240 2540 -2200
rect 2440 -2300 2460 -2240
rect 2520 -2300 2540 -2240
rect 2440 -2660 2540 -2620
rect 2440 -2720 2460 -2660
rect 2520 -2720 2540 -2660
rect 2440 -2740 2540 -2720
rect 2440 -3060 2540 -3040
rect 2440 -3120 2460 -3060
rect 2520 -3120 2540 -3060
rect 2440 -3140 2540 -3120
rect 2440 -3500 2540 -3460
rect 2440 -3560 2460 -3500
rect 2520 -3560 2540 -3500
rect 2440 -3580 2540 -3560
rect 2440 -3900 2540 -3880
rect 2440 -3960 2460 -3900
rect 2520 -3960 2540 -3900
rect 2440 -3980 2540 -3960
rect 2440 -4320 2540 -4280
rect 2440 -4380 2460 -4320
rect 2520 -4380 2540 -4320
rect 2440 -4400 2540 -4380
rect 2620 -4800 2740 -1460
rect 2840 -4500 2960 -1460
rect 3040 -1820 3142 -1800
rect 3040 -1880 3060 -1820
rect 3120 -1880 3142 -1820
rect 3040 -1900 3142 -1880
rect 3040 -2220 3140 -2200
rect 3040 -2240 3142 -2220
rect 3040 -2300 3060 -2240
rect 3120 -2300 3142 -2240
rect 3040 -2320 3142 -2300
rect 3040 -2660 3142 -2638
rect 3040 -2720 3060 -2660
rect 3120 -2720 3142 -2660
rect 3040 -2738 3142 -2720
rect 3040 -2740 3140 -2738
rect 3040 -3060 3142 -3040
rect 3040 -3120 3060 -3060
rect 3120 -3120 3142 -3060
rect 3040 -3140 3142 -3120
rect 3040 -3500 3142 -3480
rect 3040 -3560 3060 -3500
rect 3120 -3560 3142 -3500
rect 3040 -3580 3142 -3560
rect 3038 -3900 3140 -3880
rect 3038 -3960 3060 -3900
rect 3120 -3960 3140 -3900
rect 3038 -3980 3140 -3960
rect 3040 -4320 3142 -4300
rect 3040 -4380 3060 -4320
rect 3120 -4380 3142 -4320
rect 3040 -4400 3142 -4380
rect 2840 -4520 2980 -4500
rect 2840 -4580 2860 -4520
rect 2960 -4580 2980 -4520
rect 2840 -4600 2980 -4580
rect 3220 -4800 3340 -1460
rect 2020 -4840 3340 -4800
rect -420 -5060 -220 -4920
rect 2020 -4980 2820 -4840
rect 2920 -4980 3340 -4840
rect 2020 -5060 3340 -4980
<< via1 >>
rect 1860 -1440 1920 -1380
rect 500 -2220 560 -2160
rect 240 -3060 300 -3000
rect 1360 -3060 1420 -3000
rect 1860 -1880 1920 -1820
rect 1860 -2300 1920 -2240
rect 1860 -2720 1920 -2660
rect 1860 -3120 1920 -3060
rect 1860 -3560 1920 -3500
rect 1860 -3960 1920 -3900
rect 1860 -4380 1920 -4320
rect 1240 -4720 1320 -4620
rect 2460 -1440 2520 -1380
rect 3060 -1440 3120 -1380
rect 2460 -1880 2520 -1820
rect 2460 -2300 2520 -2240
rect 2460 -2720 2520 -2660
rect 2460 -3120 2520 -3060
rect 2460 -3560 2520 -3500
rect 2460 -3960 2520 -3900
rect 2460 -4380 2520 -4320
rect 3060 -1880 3120 -1820
rect 3060 -2300 3120 -2240
rect 3060 -2720 3120 -2660
rect 3060 -3120 3120 -3060
rect 3060 -3560 3120 -3500
rect 3060 -3960 3120 -3900
rect 3060 -4380 3120 -4320
rect 2860 -4580 2960 -4520
<< metal2 >>
rect 1840 -1380 1940 -1360
rect 1840 -1440 1860 -1380
rect 1920 -1440 1940 -1380
rect 1840 -1820 1940 -1440
rect 1840 -1880 1860 -1820
rect 1920 -1880 1940 -1820
rect 480 -2160 640 -2140
rect 480 -2220 500 -2160
rect 560 -2220 640 -2160
rect 480 -2660 640 -2220
rect 220 -2800 640 -2660
rect 1840 -2240 1940 -1880
rect 1840 -2300 1860 -2240
rect 1920 -2300 1940 -2240
rect 1840 -2660 1940 -2300
rect 1840 -2720 1860 -2660
rect 1920 -2720 1940 -2660
rect 220 -3000 340 -2800
rect 1840 -2980 1940 -2720
rect 220 -3060 240 -3000
rect 300 -3060 340 -3000
rect 220 -3080 340 -3060
rect 1340 -3000 1940 -2980
rect 1340 -3060 1360 -3000
rect 1420 -3060 1940 -3000
rect 1340 -3080 1860 -3060
rect 1840 -3120 1860 -3080
rect 1920 -3120 1940 -3060
rect 1840 -3500 1940 -3120
rect 1840 -3560 1860 -3500
rect 1920 -3560 1940 -3500
rect 1840 -3900 1940 -3560
rect 1840 -3960 1860 -3900
rect 1920 -3960 1940 -3900
rect 1840 -4320 1940 -3960
rect 1840 -4380 1860 -4320
rect 1920 -4380 1940 -4320
rect 1840 -4400 1940 -4380
rect 2440 -1380 2540 -1360
rect 2440 -1440 2460 -1380
rect 2520 -1440 2540 -1380
rect 2440 -1820 2540 -1440
rect 2440 -1880 2460 -1820
rect 2520 -1880 2540 -1820
rect 2440 -2240 2540 -1880
rect 2440 -2300 2460 -2240
rect 2520 -2300 2540 -2240
rect 2440 -2660 2540 -2300
rect 2440 -2720 2460 -2660
rect 2520 -2720 2540 -2660
rect 2440 -3060 2540 -2720
rect 2440 -3120 2460 -3060
rect 2520 -3120 2540 -3060
rect 2440 -3500 2540 -3120
rect 2440 -3560 2460 -3500
rect 2520 -3560 2540 -3500
rect 2440 -3900 2540 -3560
rect 3040 -1380 3140 -1360
rect 3040 -1440 3060 -1380
rect 3120 -1440 3140 -1380
rect 3040 -1820 3140 -1440
rect 3040 -1880 3060 -1820
rect 3120 -1880 3140 -1820
rect 3040 -2220 3140 -1880
rect 3040 -2240 3142 -2220
rect 3040 -2300 3060 -2240
rect 3120 -2300 3142 -2240
rect 3040 -2320 3142 -2300
rect 3040 -2638 3140 -2320
rect 3040 -2660 3142 -2638
rect 3040 -2720 3060 -2660
rect 3120 -2720 3142 -2660
rect 3040 -2738 3142 -2720
rect 3040 -3040 3140 -2738
rect 3040 -3060 3142 -3040
rect 3040 -3120 3060 -3060
rect 3120 -3120 3142 -3060
rect 3040 -3140 3142 -3120
rect 3040 -3480 3140 -3140
rect 3040 -3500 3142 -3480
rect 3040 -3560 3060 -3500
rect 3120 -3560 3142 -3500
rect 3040 -3580 3142 -3560
rect 3040 -3880 3140 -3580
rect 2440 -3960 2460 -3900
rect 2520 -3960 2540 -3900
rect 2440 -4320 2540 -3960
rect 3038 -3900 3140 -3880
rect 3038 -3960 3060 -3900
rect 3120 -3960 3140 -3900
rect 3038 -3980 3140 -3960
rect 2440 -4380 2460 -4320
rect 2520 -4380 2540 -4320
rect 2440 -4400 2540 -4380
rect 3040 -4300 3140 -3980
rect 3040 -4320 3142 -4300
rect 3040 -4380 3060 -4320
rect 3120 -4380 3142 -4320
rect 3040 -4400 3142 -4380
rect 2840 -4520 2980 -4500
rect 2840 -4580 2860 -4520
rect 2960 -4580 2980 -4520
rect 2840 -4620 2980 -4580
rect 1180 -4720 1240 -4620
rect 1320 -4720 2980 -4620
rect 1180 -4740 2980 -4720
use sky130_fd_pr__nfet_01v8_S7RYHB  XN1
timestamp 1656710231
transform 1 0 1896 0 1 -3027
box -296 -1773 296 1773
use sky130_fd_pr__nfet_01v8_S7RYHB  XN2
timestamp 1656710231
transform 1 0 2496 0 1 -3027
box -296 -1773 296 1773
use sky130_fd_pr__pfet_01v8_G8P5KT  XP1
timestamp 1656710231
transform 1 0 1296 0 1 -1881
box -296 -619 296 619
use sky130_fd_pr__pfet_01v8_G8P52V  XP2
timestamp 1656710231
transform 1 0 396 0 1 -3781
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_G8PMZT  XP3
timestamp 1656710231
transform 1 0 416 0 1 -2061
box -296 -419 296 419
use sky130_fd_pr__pfet_01v8_GYGCLT  XP4
timestamp 1656710231
transform 1 0 -864 0 1 -2041
box -696 -419 696 419
use sky130_fd_pr__nfet_01v8_S7RYHB  sky130_fd_pr__nfet_01v8_S7RYHB_0
timestamp 1656710231
transform 1 0 3096 0 1 -3027
box -296 -1773 296 1773
use sky130_fd_pr__pfet_01v8_G8P52V  sky130_fd_pr__pfet_01v8_G8P52V_0
timestamp 1656710231
transform 1 0 1276 0 1 -3781
box -296 -1019 296 1019
use sky130_fd_pr__pfet_01v8_LFNPUG  sky130_fd_pr__pfet_01v8_LFNPUG_0
timestamp 1656710231
transform 1 0 -2184 0 1 -2981
box -296 -1819 296 1819
<< labels >>
flabel metal2 520 -2600 520 -2600 0 FreeSans 800 0 0 0 d
flabel metal1 840 -3740 840 -3740 0 FreeSans 800 0 0 0 c
flabel metal1 -420 -5060 -220 -4860 0 FreeSans 1600 0 0 0 vtd
port 2 nsew
flabel metal1 -1840 -1140 -1640 -940 0 FreeSans 1600 0 0 0 vts
port 1 nsew
flabel metal1 2560 -5060 2760 -4860 0 FreeSans 1600 0 0 0 gnd
port 3 nsew
flabel metal1 -240 -1140 -40 -940 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 1588 -1414 1588 -1414 0 FreeSans 800 0 0 0 a
flabel metal1 2195 -1370 2195 -1370 0 FreeSans 800 0 0 0 b
<< end >>
