magic
tech sky130A
magscale 1 2
timestamp 1669420244
<< pwell >>
rect -616 -1198 616 1198
<< psubdiff >>
rect -580 1128 -484 1162
rect 484 1128 580 1162
rect -580 1066 -546 1128
rect 546 1066 580 1128
rect -580 -1128 -546 -1066
rect 546 -1128 580 -1066
rect -580 -1162 -484 -1128
rect 484 -1162 580 -1128
<< psubdiffcont >>
rect -484 1128 484 1162
rect -580 -1066 -546 1066
rect 546 -1066 580 1066
rect -484 -1162 484 -1128
<< xpolycontact >>
rect -450 600 -380 1032
rect -450 -1032 -380 -600
rect -284 600 -214 1032
rect -284 -1032 -214 -600
rect -118 600 -48 1032
rect -118 -1032 -48 -600
rect 48 600 118 1032
rect 48 -1032 118 -600
rect 214 600 284 1032
rect 214 -1032 284 -600
rect 380 600 450 1032
rect 380 -1032 450 -600
<< xpolyres >>
rect -450 -600 -380 600
rect -284 -600 -214 600
rect -118 -600 -48 600
rect 48 -600 118 600
rect 214 -600 284 600
rect 380 -600 450 600
<< locali >>
rect -580 1128 -484 1162
rect 484 1128 580 1162
rect -580 1066 -546 1128
rect 546 1066 580 1128
rect -580 -1128 -546 -1066
rect 546 -1128 580 -1066
rect -580 -1162 -484 -1128
rect 484 -1162 580 -1128
<< viali >>
rect -434 617 -396 1014
rect -268 617 -230 1014
rect -102 617 -64 1014
rect 64 617 102 1014
rect 230 617 268 1014
rect 396 617 434 1014
rect -434 -1014 -396 -617
rect -268 -1014 -230 -617
rect -102 -1014 -64 -617
rect 64 -1014 102 -617
rect 230 -1014 268 -617
rect 396 -1014 434 -617
<< metal1 >>
rect -440 1014 -390 1026
rect -440 617 -434 1014
rect -396 617 -390 1014
rect -440 605 -390 617
rect -274 1014 -224 1026
rect -274 617 -268 1014
rect -230 617 -224 1014
rect -274 605 -224 617
rect -108 1014 -58 1026
rect -108 617 -102 1014
rect -64 617 -58 1014
rect -108 605 -58 617
rect 58 1014 108 1026
rect 58 617 64 1014
rect 102 617 108 1014
rect 58 605 108 617
rect 224 1014 274 1026
rect 224 617 230 1014
rect 268 617 274 1014
rect 224 605 274 617
rect 390 1014 440 1026
rect 390 617 396 1014
rect 434 617 440 1014
rect 390 605 440 617
rect -440 -617 -390 -605
rect -440 -1014 -434 -617
rect -396 -1014 -390 -617
rect -440 -1026 -390 -1014
rect -274 -617 -224 -605
rect -274 -1014 -268 -617
rect -230 -1014 -224 -617
rect -274 -1026 -224 -1014
rect -108 -617 -58 -605
rect -108 -1014 -102 -617
rect -64 -1014 -58 -617
rect -108 -1026 -58 -1014
rect 58 -617 108 -605
rect 58 -1014 64 -617
rect 102 -1014 108 -617
rect 58 -1026 108 -1014
rect 224 -617 274 -605
rect 224 -1014 230 -617
rect 268 -1014 274 -617
rect 224 -1026 274 -1014
rect 390 -617 440 -605
rect 390 -1014 396 -617
rect 434 -1014 440 -617
rect 390 -1026 440 -1014
<< res0p35 >>
rect -452 -602 -378 602
rect -286 -602 -212 602
rect -120 -602 -46 602
rect 46 -602 120 602
rect 212 -602 286 602
rect 378 -602 452 602
<< properties >>
string FIXED_BBOX -563 -1145 563 1145
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 6.0 m 1 nx 6 wmin 0.350 lmin 0.50 rho 2000 val 35.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
