magic
tech sky130A
magscale 1 2
timestamp 1644769631
<< metal4 >>
rect -2509 7349 2509 7390
rect -2509 2571 2253 7349
rect 2489 2571 2509 7349
rect -2509 2530 2509 2571
rect -2509 2389 2509 2430
rect -2509 -2389 2253 2389
rect 2489 -2389 2509 2389
rect -2509 -2430 2509 -2389
rect -2509 -2571 2509 -2530
rect -2509 -7349 2253 -2571
rect 2489 -7349 2509 -2571
rect -2509 -7390 2509 -7349
<< via4 >>
rect 2253 2571 2489 7349
rect 2253 -2389 2489 2389
rect 2253 -7349 2489 -2571
<< mimcap2 >>
rect -2409 7250 2251 7290
rect -2409 2670 -1911 7250
rect 1753 2670 2251 7250
rect -2409 2630 2251 2670
rect -2409 2290 2251 2330
rect -2409 -2290 -1911 2290
rect 1753 -2290 2251 2290
rect -2409 -2330 2251 -2290
rect -2409 -2670 2251 -2630
rect -2409 -7250 -1911 -2670
rect 1753 -7250 2251 -2670
rect -2409 -7290 2251 -7250
<< mimcap2contact >>
rect -1911 2670 1753 7250
rect -1911 -2290 1753 2290
rect -1911 -7250 1753 -2670
<< metal5 >>
rect -239 7274 81 7440
rect 2211 7349 2531 7440
rect -1935 7250 1777 7274
rect -1935 2670 -1911 7250
rect 1753 2670 1777 7250
rect -1935 2646 1777 2670
rect -239 2314 81 2646
rect 2211 2571 2253 7349
rect 2489 2571 2531 7349
rect 2211 2389 2531 2571
rect -1935 2290 1777 2314
rect -1935 -2290 -1911 2290
rect 1753 -2290 1777 2290
rect -1935 -2314 1777 -2290
rect -239 -2646 81 -2314
rect 2211 -2389 2253 2389
rect 2489 -2389 2531 2389
rect 2211 -2571 2531 -2389
rect -1935 -2670 1777 -2646
rect -1935 -7250 -1911 -2670
rect 1753 -7250 1777 -2670
rect -1935 -7274 1777 -7250
rect -239 -7440 81 -7274
rect 2211 -7349 2253 -2571
rect 2489 -7349 2531 -2571
rect 2211 -7440 2531 -7349
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2509 2530 2351 7390
string parameters w 23.3 l 23.3 val 1.103k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
