** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/nmos_tb-dc.sch
**.subckt nmos_tb-dc
Va in GND 1.8
V2 out GND 3.3
XM1 out in GND GND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=7 m=7
**** begin user architecture code

.dc V2 0V 10 0.01V
.control
run
let zout= out/(-i(v2))
let id=-I(v2)
plot id
plot real(zout)
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
