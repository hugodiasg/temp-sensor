magic
tech sky130A
magscale 1 2
timestamp 1644763882
<< metal4 >>
rect -2489 7289 2489 7330
rect -2489 2551 2233 7289
rect 2469 2551 2489 7289
rect -2489 2510 2489 2551
rect -2489 2369 2489 2410
rect -2489 -2369 2233 2369
rect 2469 -2369 2489 2369
rect -2489 -2410 2489 -2369
rect -2489 -2551 2489 -2510
rect -2489 -7289 2233 -2551
rect 2469 -7289 2489 -2551
rect -2489 -7330 2489 -7289
<< via4 >>
rect 2233 2551 2469 7289
rect 2233 -2369 2469 2369
rect 2233 -7289 2469 -2551
<< mimcap2 >>
rect -2389 7190 2231 7230
rect -2389 2650 -1895 7190
rect 1737 2650 2231 7190
rect -2389 2610 2231 2650
rect -2389 2270 2231 2310
rect -2389 -2270 -1895 2270
rect 1737 -2270 2231 2270
rect -2389 -2310 2231 -2270
rect -2389 -2650 2231 -2610
rect -2389 -7190 -1895 -2650
rect 1737 -7190 2231 -2650
rect -2389 -7230 2231 -7190
<< mimcap2contact >>
rect -1895 2650 1737 7190
rect -1895 -2270 1737 2270
rect -1895 -7190 1737 -2650
<< metal5 >>
rect -239 7214 81 7380
rect 2191 7289 2511 7380
rect -1919 7190 1761 7214
rect -1919 2650 -1895 7190
rect 1737 2650 1761 7190
rect -1919 2626 1761 2650
rect -239 2294 81 2626
rect 2191 2551 2233 7289
rect 2469 2551 2511 7289
rect 2191 2369 2511 2551
rect -1919 2270 1761 2294
rect -1919 -2270 -1895 2270
rect 1737 -2270 1761 2270
rect -1919 -2294 1761 -2270
rect -239 -2626 81 -2294
rect 2191 -2369 2233 2369
rect 2469 -2369 2511 2369
rect 2191 -2551 2511 -2369
rect -1919 -2650 1761 -2626
rect -1919 -7190 -1895 -2650
rect 1737 -7190 1761 -2650
rect -1919 -7214 1761 -7190
rect -239 -7380 81 -7214
rect 2191 -7289 2233 -2551
rect 2469 -7289 2511 -2551
rect 2191 -7380 2511 -7289
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2489 2510 2331 7330
string parameters w 23.1 l 23.1 val 1.084k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
