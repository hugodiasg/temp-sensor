magic
tech sky130A
timestamp 1675570359
<< metal4 >>
rect 25859 25300 26645 25340
rect 25859 24600 25900 25300
rect 26600 24600 26645 25300
rect 25859 20815 26645 24600
<< via4 >>
rect 25900 24600 26600 25300
<< metal5 >>
rect 21600 28815 29600 29600
rect 21600 27829 28615 28615
rect 21600 22384 22384 27829
rect 22585 26845 27629 27629
rect 22585 23370 23370 26845
rect 23570 25859 26645 26645
rect 23570 24354 24354 25859
rect 25859 25300 26645 25859
rect 25859 24600 25900 25300
rect 26600 24600 26645 25300
rect 25859 24554 26645 24600
rect 26845 24354 27629 26845
rect 23570 23570 27629 24354
rect 27829 23370 28615 27829
rect 22585 22585 28615 23370
rect 28815 22384 29600 28815
rect 21600 21600 29600 22384
<< end >>
