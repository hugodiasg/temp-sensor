magic
tech sky130A
magscale 1 2
timestamp 1644161670
<< error_p >>
rect 1907 2716 2015 7484
rect 1907 -2384 2015 2384
rect 1907 -7484 2015 -2716
rect 2227 -7650 2335 7650
rect 2547 2599 2655 2821
rect 2547 2279 2655 2501
rect 2547 -2501 2655 -2279
rect 2547 -2821 2655 -2599
<< metal4 >>
rect -2633 7559 2633 7600
rect -2633 2641 2377 7559
rect 2613 2641 2633 7559
rect -2633 2600 2633 2641
rect -2633 2459 2633 2500
rect -2633 -2459 2377 2459
rect 2613 -2459 2633 2459
rect -2633 -2500 2633 -2459
rect -2633 -2641 2633 -2600
rect -2633 -7559 2377 -2641
rect 2613 -7559 2633 -2641
rect -2633 -7600 2633 -7559
<< via4 >>
rect 2377 2641 2613 7559
rect 2377 -2459 2613 2459
rect 2377 -7559 2613 -2641
<< mimcap2 >>
rect -2533 7460 2267 7500
rect -2533 2740 -2257 7460
rect 1991 2740 2267 7460
rect -2533 2700 2267 2740
rect -2533 2360 2267 2400
rect -2533 -2360 -2257 2360
rect 1991 -2360 2267 2360
rect -2533 -2400 2267 -2360
rect -2533 -2740 2267 -2700
rect -2533 -7460 -2257 -2740
rect 1991 -7460 2267 -2740
rect -2533 -7500 2267 -7460
<< mimcap2contact >>
rect -2257 2740 1991 7460
rect -2257 -2360 1991 2360
rect -2257 -7460 1991 -2740
<< metal5 >>
rect -293 7484 27 7650
rect 2227 7601 2547 7650
rect 2227 7559 2655 7601
rect -2281 7460 2015 7484
rect -2281 2740 -2257 7460
rect 1991 2740 2015 7460
rect -2281 2716 2015 2740
rect -293 2384 27 2716
rect 2227 2641 2377 7559
rect 2613 2641 2655 7559
rect 2227 2599 2655 2641
rect 2227 2501 2547 2599
rect 2227 2459 2655 2501
rect -2281 2360 2015 2384
rect -2281 -2360 -2257 2360
rect 1991 -2360 2015 2360
rect -2281 -2384 2015 -2360
rect -293 -2716 27 -2384
rect 2227 -2459 2377 2459
rect 2613 -2459 2655 2459
rect 2227 -2501 2655 -2459
rect 2227 -2599 2547 -2501
rect 2227 -2641 2655 -2599
rect -2281 -2740 2015 -2716
rect -2281 -7460 -2257 -2740
rect 1991 -7460 2015 -2740
rect -2281 -7484 2015 -7460
rect -293 -7650 27 -7484
rect 2227 -7559 2377 -2641
rect 2613 -7559 2655 -2641
rect 2227 -7601 2655 -7559
rect 2227 -7650 2547 -7601
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2633 2600 2367 7600
string parameters w 24.0 l 24.0 val 1.17k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 90
string library sky130
<< end >>
