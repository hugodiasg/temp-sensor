magic
tech sky130A
magscale 1 2
timestamp 1645495691
<< error_p >>
rect 2189 -23454 2485 23454
rect 2509 18513 2805 23405
rect 2509 18291 2829 18513
rect 2509 17971 2829 18193
rect 2509 13301 2805 17971
rect 2509 13079 2829 13301
rect 2509 12759 2829 12981
rect 2509 8089 2805 12759
rect 2509 7867 2829 8089
rect 2509 7547 2829 7769
rect 2509 2877 2805 7547
rect 2509 2655 2829 2877
rect 2509 2335 2829 2557
rect 2509 -2335 2805 2335
rect 2509 -2557 2829 -2335
rect 2509 -2877 2829 -2655
rect 2509 -7547 2805 -2877
rect 2509 -7769 2829 -7547
rect 2509 -8089 2829 -7867
rect 2509 -12759 2805 -8089
rect 2509 -12981 2829 -12759
rect 2509 -13301 2829 -13079
rect 2509 -17971 2805 -13301
rect 2509 -18193 2829 -17971
rect 2509 -18513 2829 -18291
rect 2509 -23405 2805 -18513
<< metal4 >>
rect -2807 23363 2807 23404
rect -2807 18333 2551 23363
rect 2787 18333 2807 23363
rect -2807 18292 2807 18333
rect -2807 18151 2807 18192
rect -2807 13121 2551 18151
rect 2787 13121 2807 18151
rect -2807 13080 2807 13121
rect -2807 12939 2807 12980
rect -2807 7909 2551 12939
rect 2787 7909 2807 12939
rect -2807 7868 2807 7909
rect -2807 7727 2807 7768
rect -2807 2697 2551 7727
rect 2787 2697 2807 7727
rect -2807 2656 2807 2697
rect -2807 2515 2807 2556
rect -2807 -2515 2551 2515
rect 2787 -2515 2807 2515
rect -2807 -2556 2807 -2515
rect -2807 -2697 2807 -2656
rect -2807 -7727 2551 -2697
rect 2787 -7727 2807 -2697
rect -2807 -7768 2807 -7727
rect -2807 -7909 2807 -7868
rect -2807 -12939 2551 -7909
rect 2787 -12939 2807 -7909
rect -2807 -12980 2807 -12939
rect -2807 -13121 2807 -13080
rect -2807 -18151 2551 -13121
rect 2787 -18151 2807 -13121
rect -2807 -18192 2807 -18151
rect -2807 -18333 2807 -18292
rect -2807 -23363 2551 -18333
rect 2787 -23363 2807 -18333
rect -2807 -23404 2807 -23363
<< via4 >>
rect 2551 18333 2787 23363
rect 2551 13121 2787 18151
rect 2551 7909 2787 12939
rect 2551 2697 2787 7727
rect 2551 -2515 2787 2515
rect 2551 -7727 2787 -2697
rect 2551 -12939 2787 -7909
rect 2551 -18151 2787 -13121
rect 2551 -23363 2787 -18333
<< mimcap2 >>
rect -2707 23264 2205 23304
rect -2707 18432 -2667 23264
rect 2165 18432 2205 23264
rect -2707 18392 2205 18432
rect -2707 18052 2205 18092
rect -2707 13220 -2667 18052
rect 2165 13220 2205 18052
rect -2707 13180 2205 13220
rect -2707 12840 2205 12880
rect -2707 8008 -2667 12840
rect 2165 8008 2205 12840
rect -2707 7968 2205 8008
rect -2707 7628 2205 7668
rect -2707 2796 -2667 7628
rect 2165 2796 2205 7628
rect -2707 2756 2205 2796
rect -2707 2416 2205 2456
rect -2707 -2416 -2667 2416
rect 2165 -2416 2205 2416
rect -2707 -2456 2205 -2416
rect -2707 -2796 2205 -2756
rect -2707 -7628 -2667 -2796
rect 2165 -7628 2205 -2796
rect -2707 -7668 2205 -7628
rect -2707 -8008 2205 -7968
rect -2707 -12840 -2667 -8008
rect 2165 -12840 2205 -8008
rect -2707 -12880 2205 -12840
rect -2707 -13220 2205 -13180
rect -2707 -18052 -2667 -13220
rect 2165 -18052 2205 -13220
rect -2707 -18092 2205 -18052
rect -2707 -18432 2205 -18392
rect -2707 -23264 -2667 -18432
rect 2165 -23264 2205 -18432
rect -2707 -23304 2205 -23264
<< mimcap2contact >>
rect -2667 18432 2165 23264
rect -2667 13220 2165 18052
rect -2667 8008 2165 12840
rect -2667 2796 2165 7628
rect -2667 -2416 2165 2416
rect -2667 -7628 2165 -2796
rect -2667 -12840 2165 -8008
rect -2667 -18052 2165 -13220
rect -2667 -23264 2165 -18432
<< metal5 >>
rect -411 23288 -91 23454
rect 2165 23288 2485 23454
rect -2691 23264 2485 23288
rect -2691 18432 -2667 23264
rect 2165 18432 2485 23264
rect -2691 18408 2485 18432
rect -411 18076 -91 18408
rect 2165 18076 2485 18408
rect 2509 23363 2829 23405
rect 2509 18333 2551 23363
rect 2787 18333 2829 23363
rect 2509 18291 2829 18333
rect -2691 18052 2485 18076
rect -2691 13220 -2667 18052
rect 2165 13220 2485 18052
rect -2691 13196 2485 13220
rect -411 12864 -91 13196
rect 2165 12864 2485 13196
rect 2509 18151 2829 18193
rect 2509 13121 2551 18151
rect 2787 13121 2829 18151
rect 2509 13079 2829 13121
rect -2691 12840 2485 12864
rect -2691 8008 -2667 12840
rect 2165 8008 2485 12840
rect -2691 7984 2485 8008
rect -411 7652 -91 7984
rect 2165 7652 2485 7984
rect 2509 12939 2829 12981
rect 2509 7909 2551 12939
rect 2787 7909 2829 12939
rect 2509 7867 2829 7909
rect -2691 7628 2485 7652
rect -2691 2796 -2667 7628
rect 2165 2796 2485 7628
rect -2691 2772 2485 2796
rect -411 2440 -91 2772
rect 2165 2440 2485 2772
rect 2509 7727 2829 7769
rect 2509 2697 2551 7727
rect 2787 2697 2829 7727
rect 2509 2655 2829 2697
rect -2691 2416 2485 2440
rect -2691 -2416 -2667 2416
rect 2165 -2416 2485 2416
rect -2691 -2440 2485 -2416
rect -411 -2772 -91 -2440
rect 2165 -2772 2485 -2440
rect 2509 2515 2829 2557
rect 2509 -2515 2551 2515
rect 2787 -2515 2829 2515
rect 2509 -2557 2829 -2515
rect -2691 -2796 2485 -2772
rect -2691 -7628 -2667 -2796
rect 2165 -7628 2485 -2796
rect -2691 -7652 2485 -7628
rect -411 -7984 -91 -7652
rect 2165 -7984 2485 -7652
rect 2509 -2697 2829 -2655
rect 2509 -7727 2551 -2697
rect 2787 -7727 2829 -2697
rect 2509 -7769 2829 -7727
rect -2691 -8008 2485 -7984
rect -2691 -12840 -2667 -8008
rect 2165 -12840 2485 -8008
rect -2691 -12864 2485 -12840
rect -411 -13196 -91 -12864
rect 2165 -13196 2485 -12864
rect 2509 -7909 2829 -7867
rect 2509 -12939 2551 -7909
rect 2787 -12939 2829 -7909
rect 2509 -12981 2829 -12939
rect -2691 -13220 2485 -13196
rect -2691 -18052 -2667 -13220
rect 2165 -18052 2485 -13220
rect -2691 -18076 2485 -18052
rect -411 -18408 -91 -18076
rect 2165 -18408 2485 -18076
rect 2509 -13121 2829 -13079
rect 2509 -18151 2551 -13121
rect 2787 -18151 2829 -13121
rect 2509 -18193 2829 -18151
rect -2691 -18432 2485 -18408
rect -2691 -23264 -2667 -18432
rect 2165 -23264 2485 -18432
rect -2691 -23288 2485 -23264
rect -411 -23454 -91 -23288
rect 2165 -23454 2485 -23288
rect 2509 -18333 2829 -18291
rect 2509 -23363 2551 -18333
rect 2787 -23363 2829 -18333
rect 2509 -23405 2829 -23363
<< properties >>
string FIXED_BBOX -2807 18292 2305 23404
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.559 l 24.559 val 1.224k carea 2.00 cperi 0.19 nx 1 ny 9 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
