magic
tech sky130A
magscale 1 2
timestamp 1645800166
<< metal4 >>
rect -2622 7688 2622 7729
rect -2622 2684 2366 7688
rect 2602 2684 2622 7688
rect -2622 2643 2622 2684
rect -2622 2502 2622 2543
rect -2622 -2502 2366 2502
rect 2602 -2502 2622 2502
rect -2622 -2543 2622 -2502
rect -2622 -2684 2622 -2643
rect -2622 -7688 2366 -2684
rect 2602 -7688 2622 -2684
rect -2622 -7729 2622 -7688
<< via4 >>
rect 2366 2684 2602 7688
rect 2366 -2502 2602 2502
rect 2366 -7688 2602 -2684
<< mimcap2 >>
rect -2522 7589 2364 7629
rect -2522 2783 -2001 7589
rect 1843 2783 2364 7589
rect -2522 2743 2364 2783
rect -2522 2403 2364 2443
rect -2522 -2403 -2001 2403
rect 1843 -2403 2364 2403
rect -2522 -2443 2364 -2403
rect -2522 -2783 2364 -2743
rect -2522 -7589 -2001 -2783
rect 1843 -7589 2364 -2783
rect -2522 -7629 2364 -7589
<< mimcap2contact >>
rect -2001 2783 1843 7589
rect -2001 -2403 1843 2403
rect -2001 -7589 1843 -2783
<< metal5 >>
rect -239 7613 81 7779
rect 2324 7688 2644 7779
rect -2025 7589 1867 7613
rect -2025 2783 -2001 7589
rect 1843 2783 1867 7589
rect -2025 2759 1867 2783
rect -239 2427 81 2759
rect 2324 2684 2366 7688
rect 2602 2684 2644 7688
rect 2324 2502 2644 2684
rect -2025 2403 1867 2427
rect -2025 -2403 -2001 2403
rect 1843 -2403 1867 2403
rect -2025 -2427 1867 -2403
rect -239 -2759 81 -2427
rect 2324 -2502 2366 2502
rect 2602 -2502 2644 2502
rect 2324 -2684 2644 -2502
rect -2025 -2783 1867 -2759
rect -2025 -7589 -2001 -2783
rect 1843 -7589 1867 -2783
rect -2025 -7613 1867 -7589
rect -239 -7779 81 -7613
rect 2324 -7688 2366 -2684
rect 2602 -7688 2644 -2684
rect 2324 -7779 2644 -7688
<< properties >>
string FIXED_BBOX -2622 2643 2464 7729
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.43 l 24.43 val 1.212k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
