magic
tech sky130A
magscale 1 2
timestamp 1669916246
<< pwell >>
rect -296 -310 296 310
<< nmos >>
rect -100 -100 100 100
<< ndiff >>
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
<< ndiffc >>
rect -146 -88 -112 88
rect 112 -88 146 88
<< psubdiff >>
rect -260 240 -164 274
rect 164 240 260 274
rect -260 178 -226 240
rect 226 178 260 240
rect -260 -240 -226 -178
rect 226 -240 260 -178
rect -260 -274 -164 -240
rect 164 -274 260 -240
<< psubdiffcont >>
rect -164 240 164 274
rect -260 -178 -226 178
rect 226 -178 260 178
rect -164 -274 164 -240
<< poly >>
rect -100 172 100 188
rect -100 138 -84 172
rect 84 138 100 172
rect -100 100 100 138
rect -100 -138 100 -100
rect -100 -172 -84 -138
rect 84 -172 100 -138
rect -100 -188 100 -172
<< polycont >>
rect -84 138 84 172
rect -84 -172 84 -138
<< locali >>
rect -260 240 -164 274
rect 164 240 260 274
rect -260 178 -226 240
rect 226 178 260 240
rect -100 138 -84 172
rect 84 138 100 172
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect -100 -172 -84 -138
rect 84 -172 100 -138
rect -260 -274 -226 -178
rect 226 -274 260 -178
<< viali >>
rect -59 138 59 172
rect -146 -88 -112 88
rect 112 -88 146 88
rect -59 -172 59 -138
rect -226 -274 -164 -240
rect -164 -274 164 -240
rect 164 -274 226 -240
<< metal1 >>
rect -71 172 71 178
rect -71 138 -59 172
rect 59 138 71 172
rect -71 132 71 138
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect -71 -138 71 -132
rect -71 -172 -59 -138
rect 59 -172 71 -138
rect -71 -178 71 -172
rect -238 -240 238 -234
rect -238 -274 -226 -240
rect 226 -274 238 -240
rect -238 -280 238 -274
<< properties >>
string FIXED_BBOX -243 -257 243 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
