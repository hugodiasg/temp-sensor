magic
tech sky130A
magscale 1 2
timestamp 1700775626
<< metal1 >>
rect 6780 16240 6980 16420
rect 6780 16140 7000 16240
rect 6590 15520 6600 16140
rect 7200 15520 7210 16140
rect 6570 13880 6580 14480
rect 7180 13880 7190 14480
rect 660 -5520 860 -5460
rect 660 -5600 1660 -5520
rect 660 -5660 860 -5600
rect 1600 -5940 1660 -5600
rect 950 -6000 960 -5940
rect 660 -6200 960 -6000
rect 950 -6260 960 -6200
rect 1240 -6000 1250 -5940
rect 1240 -6200 1580 -6000
rect 1240 -6260 1250 -6200
rect 1680 -6340 1980 -6000
rect 1600 -6460 1660 -6400
rect 1780 -10360 1980 -6340
<< via1 >>
rect 6600 15520 7200 16140
rect 6580 13880 7180 14480
rect 960 -6260 1240 -5940
<< metal2 >>
rect 6600 16140 7200 16150
rect 6600 15510 7200 15520
rect 6580 14480 7180 14490
rect 6580 13870 7180 13880
rect 960 -5940 1240 -5930
rect 960 -6270 1240 -6260
<< via2 >>
rect 6600 15520 7200 16140
rect 6580 13880 7180 14480
rect 960 -6260 1240 -5940
<< metal3 >>
rect 6590 16140 7210 16145
rect 6590 15520 6600 16140
rect 7200 15520 7210 16140
rect 6590 15515 7210 15520
rect 6570 14480 7190 14485
rect 6570 13880 6580 14480
rect 7180 13880 7190 14480
rect 6570 13875 7190 13880
rect 950 -5940 1250 -5935
rect 950 -6260 960 -5940
rect 1240 -6260 1250 -5940
rect 950 -6265 1250 -6260
rect 860 -7880 23078 -7800
rect 860 -10080 900 -7880
rect 1340 -8020 23078 -7880
rect 1340 -10040 20940 -8020
rect 22860 -10040 23078 -8020
rect 1340 -10080 23078 -10040
rect 860 -10160 23078 -10080
<< via3 >>
rect 6600 15520 7200 16140
rect 6580 13880 7180 14480
rect 960 -6260 1240 -5940
rect 900 -10080 1340 -7880
rect 20940 -10040 22860 -8020
<< metal4 >>
rect 6599 16140 7201 16141
rect 6599 15520 6600 16140
rect 7200 15520 7201 16140
rect 6599 15519 7201 15520
rect 6579 14480 7181 14481
rect 6579 13880 6580 14480
rect 7180 13880 7181 14480
rect 6579 13879 7181 13880
rect 840 -5940 1380 580
rect 840 -6260 960 -5940
rect 1240 -6260 1380 -5940
rect 840 -7880 1380 -6260
rect 840 -10080 900 -7880
rect 1340 -10080 1380 -7880
rect 20939 -8020 22861 -8019
rect 20939 -10040 20940 -8020
rect 22860 -10040 22861 -8020
rect 20939 -10041 22861 -10040
rect 840 -10160 1380 -10080
<< via4 >>
rect 6600 15520 7200 16140
rect 6580 13880 7180 14480
<< metal5 >>
rect 5679 16140 9782 16202
rect 5679 15520 6600 16140
rect 7200 15520 9782 16140
rect 5679 14480 9782 15520
rect 5679 13880 6580 14480
rect 7180 13880 9782 14480
rect 5679 13840 9782 13880
<< comment >>
rect 7400 -10160 7420 -10140
use l0  l0_0
timestamp 1700108998
transform 1 0 -31780 0 1 -46998
box 39200 36838 63200 63200
use sky130_fd_pr__cap_mim_m3_2_5FNSJ7  XC0
timestamp 1700108998
transform -1 0 3651 0 -1 8320
box -2789 -7920 2811 7920
use sky130_fd_pr__nfet_01v8_LPSAWK  XM1
timestamp 1700142087
transform 1 0 1631 0 1 -6170
box -211 -410 211 410
use sky130_fd_pr__res_xhigh_po_0p35_7RFGLT  XR1
timestamp 1700108998
transform 1 0 6901 0 1 13398
box -201 -1098 201 1098
<< labels >>
flabel metal1 6780 16220 6980 16420 0 FreeSans 256 0 0 0 vd
port 3 nsew
flabel metal1 1780 -10360 1980 -10160 0 FreeSans 256 0 0 0 gnd
port 0 nsew
flabel metal1 660 -6200 860 -6000 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 660 -5660 860 -5460 0 FreeSans 256 0 0 0 in
port 1 nsew
<< end >>
