magic
tech sky130B
timestamp 1644922882
<< metal4 >>
rect -1255 3674 1254 3695
rect -1255 1285 1126 3674
rect 1244 1285 1254 3674
rect -1255 1265 1254 1285
rect -1255 1194 1254 1215
rect -1255 -1195 1126 1194
rect 1244 -1195 1254 1194
rect -1255 -1215 1254 -1195
rect -1255 -1286 1254 -1265
rect -1255 -3675 1126 -1286
rect 1244 -3675 1254 -1286
rect -1255 -3695 1254 -3675
<< via4 >>
rect 1126 1285 1244 3674
rect 1126 -1195 1244 1194
rect 1126 -3675 1244 -1286
<< mimcap2 >>
rect -1205 3625 1125 3645
rect -1205 1335 -956 3625
rect 876 1335 1125 3625
rect -1205 1315 1125 1335
rect -1205 1145 1125 1165
rect -1205 -1145 -956 1145
rect 876 -1145 1125 1145
rect -1205 -1165 1125 -1145
rect -1205 -1335 1125 -1315
rect -1205 -3625 -956 -1335
rect 876 -3625 1125 -1335
rect -1205 -3645 1125 -3625
<< mimcap2contact >>
rect -956 1335 876 3625
rect -956 -1145 876 1145
rect -956 -3625 876 -1335
<< metal5 >>
rect -120 3637 40 3720
rect 1105 3674 1265 3720
rect -968 3625 888 3637
rect -968 1335 -956 3625
rect 876 1335 888 3625
rect -968 1323 888 1335
rect -120 1157 40 1323
rect 1105 1285 1126 3674
rect 1244 1285 1265 3674
rect 1105 1194 1265 1285
rect -968 1145 888 1157
rect -968 -1145 -956 1145
rect 876 -1145 888 1145
rect -968 -1157 888 -1145
rect -120 -1323 40 -1157
rect 1105 -1195 1126 1194
rect 1244 -1195 1265 1194
rect 1105 -1286 1265 -1195
rect -968 -1335 888 -1323
rect -968 -3625 -956 -1335
rect 876 -3625 888 -1335
rect -968 -3637 888 -3625
rect -120 -3720 40 -3637
rect 1105 -3675 1126 -1286
rect 1244 -3675 1265 -1286
rect 1105 -3720 1265 -3675
<< properties >>
string FIXED_BBOX -628 632 587 1847
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.3 l 23.3 val 1.103k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
