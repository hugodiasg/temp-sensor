magic
tech sky130A
magscale 1 2
timestamp 1700764089
<< nwell >>
rect 1140 4880 7520 5620
rect 1167 2127 2533 4880
rect 6160 2120 7520 4880
<< pwell >>
rect 2840 4080 6032 4860
rect 2840 3640 4220 4080
rect 4240 3640 6032 4080
rect 2840 2660 6032 3640
<< psubdiff >>
rect 2876 4810 2972 4844
rect 5900 4810 5996 4844
rect 2876 4748 2910 4810
rect 2876 2730 2910 2792
rect 5962 4748 5996 4810
rect 5962 2730 5996 2792
rect 2876 2696 2972 2730
rect 5900 2696 5996 2730
<< nsubdiff >>
rect 7380 5577 7480 5580
rect 1203 5543 1263 5577
rect 7417 5543 7480 5577
rect 1203 5517 1237 5543
rect 2603 5540 2637 5543
rect 6103 5540 6137 5543
rect 7380 5540 7480 5543
rect 7443 5517 7477 5540
rect 2480 4957 2740 4960
rect 6203 4957 6237 4960
rect 1237 4923 1240 4957
rect 2460 4923 2680 4957
rect 6060 4923 6237 4957
rect 7440 4923 7443 4957
rect 2460 4920 2740 4923
rect 2460 4843 2497 4920
rect 6203 4880 6237 4923
rect 1203 2197 1237 2223
rect 2463 4840 2497 4843
rect 2463 2197 2497 2223
rect 1203 2163 1263 2197
rect 2437 2163 2497 2197
rect 6203 2197 6237 2223
rect 7443 2197 7477 2223
rect 6203 2163 6263 2197
rect 7417 2163 7477 2197
<< psubdiffcont >>
rect 2972 4810 5900 4844
rect 2876 2792 2910 4748
rect 5962 2792 5996 4748
rect 2972 2696 5900 2730
<< nsubdiffcont >>
rect 1263 5543 7417 5577
rect 1203 2223 1237 5517
rect 2680 4923 6060 4957
rect 2463 2223 2497 4840
rect 1263 2163 2437 2197
rect 6203 2223 6237 4880
rect 7443 2223 7477 5517
rect 6263 2163 7417 2197
<< locali >>
rect 7380 5577 7480 5580
rect 1203 5543 1263 5577
rect 7417 5543 7480 5577
rect 1203 5517 1237 5543
rect 2603 5540 2637 5543
rect 6103 5540 6137 5543
rect 7380 5540 7480 5543
rect 7443 5517 7477 5540
rect 2480 4957 2740 4960
rect 6203 4957 6237 4960
rect 1237 4923 1240 4957
rect 2460 4923 2680 4957
rect 6060 4923 6237 4957
rect 7440 4923 7443 4957
rect 2460 4920 2740 4923
rect 2460 4843 2497 4920
rect 6203 4880 6237 4923
rect 2463 4840 2497 4843
rect 1203 2197 1237 2223
rect 2876 4810 2972 4844
rect 5900 4810 5996 4844
rect 2876 4748 2910 4810
rect 2876 2730 2910 2792
rect 5962 4748 5996 4810
rect 5962 2730 5996 2792
rect 2876 2696 2972 2730
rect 5900 2696 5996 2730
rect 2463 2197 2497 2223
rect 1203 2163 1263 2197
rect 2437 2163 2497 2197
rect 6203 2197 6237 2223
rect 7443 2197 7477 2223
rect 6203 2163 6263 2197
rect 7417 2163 7477 2197
<< viali >>
rect 3820 5577 4860 5580
rect 3820 5543 4860 5577
rect 3820 5540 4860 5543
rect 1628 5407 1796 5441
rect 1886 5407 2054 5441
rect 2788 5407 2956 5441
rect 5740 5407 5908 5441
rect 6628 5407 6796 5441
rect 6886 5407 7054 5441
rect 2530 5079 2698 5113
rect 2788 5079 2956 5113
rect 3046 5079 3214 5113
rect 3304 5079 3472 5113
rect 3562 5079 3730 5113
rect 3820 5079 3988 5113
rect 4078 5079 4246 5113
rect 4470 5079 4638 5113
rect 4728 5079 4896 5113
rect 4986 5079 5154 5113
rect 5244 5079 5412 5113
rect 5502 5079 5670 5113
rect 5740 5079 5908 5113
rect 5998 5079 6186 5113
rect 1370 2279 1538 2313
rect 2144 2279 2312 2313
rect 3640 2730 3740 2760
rect 5060 2730 5160 2760
rect 3640 2696 3740 2730
rect 5060 2696 5160 2730
rect 3640 2680 3740 2696
rect 5060 2680 5160 2696
rect 6370 2279 6538 2313
rect 7144 2279 7312 2313
<< metal1 >>
rect 1800 5520 1820 5640
rect 1880 5620 4000 5640
rect 4280 5620 4480 5820
rect 1880 5520 3720 5620
rect 3820 5580 4860 5620
rect 3820 5520 4860 5540
rect 4960 5600 6900 5620
rect 4960 5520 6800 5600
rect 1800 5500 6800 5520
rect 6860 5500 6900 5600
rect 1616 5441 1808 5447
rect 1616 5440 1628 5441
rect 1360 5407 1628 5440
rect 1796 5440 1808 5441
rect 1874 5441 2066 5447
rect 1874 5440 1886 5441
rect 1796 5407 1886 5440
rect 2054 5440 2066 5441
rect 2776 5441 2968 5447
rect 2776 5440 2788 5441
rect 2054 5407 2788 5440
rect 2956 5407 2968 5441
rect 1360 5401 2968 5407
rect 5720 5441 7320 5460
rect 5720 5407 5740 5441
rect 5908 5407 6628 5441
rect 6796 5407 6886 5441
rect 7054 5407 7320 5441
rect 1360 5400 2960 5401
rect 5720 5400 7320 5407
rect 2720 5320 3720 5360
rect 1790 4960 1800 5200
rect 1900 4960 1910 5200
rect 2480 5113 2740 5320
rect 3710 5280 3720 5320
rect 3820 5280 3830 5360
rect 4040 5260 4300 5360
rect 4660 5320 5720 5360
rect 3990 5200 4000 5260
rect 2960 5160 4000 5200
rect 4080 5160 4300 5260
rect 3800 5120 4000 5160
rect 2780 5119 4000 5120
rect 2480 5080 2530 5113
rect 2518 5079 2530 5080
rect 2698 5080 2740 5113
rect 2776 5113 4000 5119
rect 2698 5079 2710 5080
rect 2518 5073 2710 5079
rect 2776 5079 2788 5113
rect 2956 5080 3046 5113
rect 2956 5079 2968 5080
rect 2776 5073 2968 5079
rect 3034 5079 3046 5080
rect 3214 5080 3304 5113
rect 3214 5079 3226 5080
rect 3034 5073 3226 5079
rect 3292 5079 3304 5080
rect 3472 5080 3562 5113
rect 3472 5079 3484 5080
rect 3292 5073 3484 5079
rect 3550 5079 3562 5080
rect 3730 5080 3820 5113
rect 3730 5079 3742 5080
rect 3550 5073 3742 5079
rect 3808 5079 3820 5080
rect 3988 5079 4000 5113
rect 4040 5113 4300 5160
rect 4040 5080 4078 5113
rect 3808 5073 4000 5079
rect 4066 5079 4078 5080
rect 4246 5080 4300 5113
rect 4420 5240 4640 5320
rect 4720 5240 4730 5320
rect 6080 5280 6240 5340
rect 4420 5180 4680 5240
rect 4420 5120 4740 5180
rect 4870 5160 4880 5280
rect 4960 5200 4970 5280
rect 5940 5240 6240 5280
rect 5940 5200 6220 5240
rect 4960 5160 6220 5200
rect 4420 5119 5900 5120
rect 4420 5113 5920 5119
rect 4420 5080 4470 5113
rect 4246 5079 4258 5080
rect 4066 5073 4258 5079
rect 4458 5079 4470 5080
rect 4638 5080 4728 5113
rect 4638 5079 4650 5080
rect 4458 5073 4650 5079
rect 4716 5079 4728 5080
rect 4896 5080 4986 5113
rect 4896 5079 4908 5080
rect 4716 5073 4908 5079
rect 4974 5079 4986 5080
rect 5154 5080 5244 5113
rect 5154 5079 5166 5080
rect 4974 5073 5166 5079
rect 5232 5079 5244 5080
rect 5412 5080 5502 5113
rect 5412 5079 5424 5080
rect 5232 5073 5424 5079
rect 5490 5079 5502 5080
rect 5670 5080 5740 5113
rect 5670 5079 5682 5080
rect 5490 5073 5682 5079
rect 5728 5079 5740 5080
rect 5908 5079 5920 5113
rect 5980 5113 6220 5160
rect 5980 5100 5998 5113
rect 5728 5073 5920 5079
rect 5986 5079 5998 5100
rect 6186 5080 6220 5113
rect 6186 5079 6198 5080
rect 5986 5073 6198 5079
rect 4290 4820 4300 4900
rect 4380 4820 6060 4900
rect 6140 4820 6150 4900
rect 4290 4720 4300 4780
rect 4380 4720 4390 4780
rect 4500 4740 4560 4780
rect 6790 4760 6800 5320
rect 6860 4760 6870 5320
rect 4480 4680 4580 4740
rect 3990 4600 4000 4680
rect 4080 4600 4280 4680
rect 4160 4400 4280 4600
rect 4480 4600 4640 4680
rect 4720 4600 4730 4680
rect 4330 4400 4340 4480
rect 4400 4400 4410 4480
rect 4480 4460 4580 4600
rect 4200 4300 4280 4400
rect 4400 4340 4460 4360
rect 4630 4340 4640 4360
rect 4400 4300 4640 4340
rect 4700 4340 4710 4360
rect 4700 4300 4720 4340
rect 2570 4180 2580 4240
rect 2640 4180 4640 4240
rect 4700 4180 4720 4240
rect 3910 4080 3920 4140
rect 4000 4080 4340 4140
rect 4400 4080 4410 4140
rect 1300 3760 1580 3940
rect 2080 3760 2360 3940
rect 3220 3900 3360 4040
rect 4000 3960 4200 4040
rect 3940 3940 4200 3960
rect 3140 3820 3440 3900
rect 3520 3820 3530 3900
rect 3220 3700 3360 3820
rect 3440 3740 3520 3820
rect 3630 3780 3640 3880
rect 3740 3780 3750 3880
rect 3910 3840 3920 3940
rect 3980 3840 4200 3940
rect 4320 3840 4540 3980
rect 4640 3940 5580 4000
rect 4640 3880 4840 3940
rect 3940 3820 4200 3840
rect 3440 3700 3920 3740
rect 4000 3700 4200 3820
rect 4640 3780 4680 3880
rect 4380 3760 4680 3780
rect 4380 3700 4400 3760
rect 4460 3700 4680 3760
rect 4740 3780 4840 3880
rect 5660 3800 5880 3980
rect 4740 3700 4860 3780
rect 6300 3740 6600 3920
rect 7060 3740 7360 3920
rect 4380 3680 4860 3700
rect 5340 3640 5800 3660
rect 5340 3580 5720 3640
rect 5780 3580 5800 3640
rect 5340 3560 5800 3580
rect 4300 3320 4600 3440
rect 5600 3380 5880 3440
rect 7560 3280 7760 3340
rect 5740 3260 6060 3280
rect 1580 3200 4470 3220
rect 5730 3200 5740 3260
rect 5800 3220 6060 3260
rect 6120 3220 7760 3280
rect 5800 3200 7760 3220
rect 1580 3140 4400 3200
rect 4460 3140 4470 3200
rect 1580 3120 4470 3140
rect 4580 3180 5620 3200
rect 4580 3100 5060 3180
rect 4360 2860 4580 3020
rect 5050 2940 5060 3100
rect 5120 3100 5620 3180
rect 7560 3140 7760 3200
rect 5120 2940 5130 3100
rect 5620 2840 5800 2980
rect 3628 2760 3752 2766
rect 3628 2680 3640 2760
rect 3740 2680 3752 2760
rect 3628 2674 3752 2680
rect 5048 2760 5172 2766
rect 5048 2680 5060 2760
rect 5160 2680 5172 2760
rect 5048 2674 5172 2680
rect 1560 2320 1620 2620
rect 2080 2320 2140 2620
rect 6560 2340 6620 2540
rect 7080 2340 7140 2540
rect 1360 2319 2320 2320
rect 6340 2319 7320 2340
rect 1358 2313 2324 2319
rect 1358 2279 1370 2313
rect 1538 2280 2144 2313
rect 1538 2279 1550 2280
rect 1358 2273 1550 2279
rect 2132 2279 2144 2280
rect 2312 2279 2324 2313
rect 6340 2313 7324 2319
rect 6340 2280 6370 2313
rect 2132 2273 2324 2279
rect 6358 2279 6370 2280
rect 6538 2280 7144 2313
rect 6538 2279 6550 2280
rect 6358 2273 6550 2279
rect 7132 2279 7144 2280
rect 7312 2279 7324 2313
rect 7132 2273 7324 2279
rect 900 2180 1100 2220
rect 900 2100 2580 2180
rect 2640 2100 2650 2180
rect 900 2020 1100 2100
rect 900 1860 1100 1900
rect 900 1740 3440 1860
rect 3520 1740 3530 1860
rect 900 1700 1100 1740
rect 900 -1580 5180 -1520
rect 900 -1640 3660 -1580
rect 3720 -1640 5080 -1580
rect 5140 -1640 5180 -1580
rect 900 -1720 5180 -1640
<< via1 >>
rect 1820 5520 1880 5640
rect 3720 5520 3820 5620
rect 4860 5520 4960 5620
rect 6800 5500 6860 5600
rect 1800 4960 1900 5200
rect 3720 5280 3820 5360
rect 4000 5160 4080 5260
rect 4640 5240 4720 5320
rect 4880 5160 4960 5280
rect 4300 4820 4380 4900
rect 6060 4820 6140 4900
rect 4300 4720 4380 4780
rect 6800 4760 6860 5320
rect 4000 4600 4080 4680
rect 4640 4600 4720 4680
rect 4340 4400 4400 4480
rect 4640 4300 4700 4360
rect 2580 4180 2640 4240
rect 4640 4180 4700 4240
rect 3920 4080 4000 4140
rect 4340 4080 4400 4140
rect 3440 3820 3520 3900
rect 3640 3780 3740 3880
rect 3920 3840 3980 3940
rect 4400 3700 4460 3760
rect 4680 3700 4740 3880
rect 5720 3580 5780 3640
rect 5740 3200 5800 3260
rect 6060 3220 6120 3280
rect 4400 3140 4460 3200
rect 5060 2940 5120 3180
rect 3640 2680 3740 2760
rect 5060 2680 5160 2760
rect 2580 2100 2640 2180
rect 3440 1740 3520 1860
rect 3660 -1640 3720 -1580
rect 5080 -1640 5140 -1580
<< metal2 >>
rect 1820 5640 1880 5650
rect 1800 5520 1820 5640
rect 1880 5520 1900 5640
rect 1800 5200 1900 5520
rect 3720 5620 3820 5630
rect 3720 5360 3820 5520
rect 4860 5620 4960 5630
rect 4640 5320 4720 5330
rect 3720 5270 3820 5280
rect 1800 4950 1900 4960
rect 4000 5260 4080 5280
rect 4000 4680 4080 5160
rect 4300 4900 4380 4910
rect 4300 4780 4380 4820
rect 4300 4710 4380 4720
rect 4000 4590 4080 4600
rect 4640 4680 4720 5240
rect 4860 5280 4960 5520
rect 4860 5160 4880 5280
rect 4880 5150 4960 5160
rect 6780 5600 6880 5620
rect 6780 5500 6800 5600
rect 6860 5500 6880 5600
rect 6780 5320 6880 5500
rect 4640 4590 4720 4600
rect 6060 4900 6140 4910
rect 4340 4480 4400 4490
rect 2580 4240 2640 4250
rect 2580 2180 2640 4180
rect 3920 4140 4000 4150
rect 3920 3940 4000 4080
rect 4340 4140 4400 4400
rect 4640 4360 4700 4370
rect 4700 4300 4720 4340
rect 4640 4240 4720 4300
rect 4700 4180 4720 4240
rect 4640 4160 4720 4180
rect 4340 4070 4400 4080
rect 2580 2090 2640 2100
rect 3440 3900 3520 3910
rect 3440 1860 3520 3820
rect 3440 1730 3520 1740
rect 3640 3880 3740 3890
rect 3980 3840 4000 3940
rect 4680 3880 4740 3890
rect 3920 3830 3980 3840
rect 3640 2760 3740 3780
rect 4380 3760 4480 3780
rect 4380 3700 4400 3760
rect 4460 3700 4480 3760
rect 4380 3200 4480 3700
rect 4380 3140 4400 3200
rect 4460 3140 4480 3200
rect 4380 3120 4480 3140
rect 4660 3700 4680 3880
rect 4740 3700 4760 3880
rect 3640 -1580 3740 2680
rect 4660 2350 4760 3700
rect 5720 3640 5780 3650
rect 5780 3580 5800 3640
rect 5720 3260 5800 3580
rect 5720 3200 5740 3260
rect 5060 3180 5160 3200
rect 5740 3190 5800 3200
rect 6060 3280 6140 4820
rect 6780 4760 6800 5320
rect 6860 4760 6880 5320
rect 6780 4720 6880 4760
rect 6120 3220 6140 3280
rect 5120 2940 5160 3180
rect 5060 2760 5160 2940
rect 4540 2340 4960 2350
rect 4540 2050 4960 2060
rect 3640 -1640 3660 -1580
rect 3720 -1640 3740 -1580
rect 3640 -1660 3740 -1640
rect 5060 -1580 5160 2680
rect 6060 2160 6140 3220
rect 5860 2140 6340 2160
rect 5860 1880 5880 2140
rect 6320 1880 6340 2140
rect 5860 1860 6340 1880
rect 5060 -1640 5080 -1580
rect 5140 -1640 5160 -1580
rect 5060 -1660 5160 -1640
<< via2 >>
rect 4540 2060 4960 2340
rect 5880 1880 6320 2140
<< metal3 >>
rect 4530 2340 4970 2345
rect 4530 2060 4540 2340
rect 4960 2060 4970 2340
rect 4530 2055 4970 2060
rect 5860 2140 6340 2160
rect 4580 2040 4860 2055
rect 5860 1880 5880 2140
rect 6320 1880 6340 2140
rect 5860 1860 6340 1880
<< via3 >>
rect 4540 2060 4960 2340
rect 5880 1880 6320 2140
<< metal4 >>
rect 4520 2340 4980 2360
rect 4520 2060 4540 2340
rect 4960 2060 4980 2340
rect 4520 1380 4980 2060
rect 5860 2140 6340 2160
rect 5860 1860 5880 2140
rect 6320 1860 6340 2140
<< via4 >>
rect 5880 1880 6320 2140
rect 5880 1780 6320 1880
<< metal5 >>
rect 5840 2140 6360 2180
rect 5840 1780 5880 2140
rect 6320 1780 6360 2140
rect 5840 1400 6360 1780
use sky130_fd_pr__cap_mim_m3_2_26U9NK  sky130_fd_pr__cap_mim_m3_2_26U9NK_0
timestamp 1700708449
transform 1 0 4249 0 1 81
box -3349 -1581 3371 1581
use sky130_fd_pr__nfet_01v8_5VPKLS  sky130_fd_pr__nfet_01v8_5VPKLS_0
timestamp 1700704221
transform 1 0 3685 0 1 3868
box -545 -188 545 188
use sky130_fd_pr__nfet_01v8_HD5U9F  sky130_fd_pr__nfet_01v8_HD5U9F_1
timestamp 1700704221
transform 1 0 4381 0 1 4538
box -221 -238 221 238
use sky130_fd_pr__pfet_01v8_99C25S  sky130_fd_pr__pfet_01v8_99C25S_0
timestamp 1700762700
transform 1 0 1841 0 1 3860
box -581 -1600 581 1600
use sky130_fd_pr__pfet_01v8_99C25S  sky130_fd_pr__pfet_01v8_99C25S_1
timestamp 1700762700
transform 1 0 6841 0 1 3860
box -581 -1600 581 1600
use sky130_fd_pr__pfet_01v8_AXJJQ9  sky130_fd_pr__pfet_01v8_AXJJQ9_0
timestamp 1700746600
transform 1 0 3388 0 1 5260
box -968 -200 968 200
use sky130_fd_pr__pfet_01v8_AXJJQ9  sky130_fd_pr__pfet_01v8_AXJJQ9_1
timestamp 1700746600
transform 1 0 5308 0 1 5260
box -968 -200 968 200
use sky130_fd_pr__nfet_01v8_MMM6UU  XM10
timestamp 1700762700
transform 1 0 5103 0 1 3408
box -803 -588 803 588
<< labels >>
flabel metal2 4020 4920 4040 4960 0 FreeSans 800 0 0 0 a
flabel metal2 4660 4920 4700 4940 0 FreeSans 800 0 0 0 b
flabel metal1 4280 5620 4480 5820 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal1 4100 4100 4120 4120 0 FreeSans 800 0 0 0 c
flabel metal1 900 1700 1100 1900 0 FreeSans 256 0 0 0 ib
port 1 nsew
flabel metal1 900 2020 1100 2220 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 2720 3180 2740 3200 0 FreeSans 800 0 0 0 d
flabel metal1 7560 3140 7760 3340 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 900 -1720 1100 -1520 0 FreeSans 256 0 0 0 gnd
port 4 nsew
<< end >>
