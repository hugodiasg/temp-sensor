** sch_path: /home/hugodg/.xschem/simulations/untitled.sch
**.subckt untitled
vpwr vpwr GND 1.8
.save i(vpwr)
V3 clk GND pulse 0 1.8 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 '
x1 vpwr clk out vts vpwr GND vd sigma-delta
vd vd GND 1.8
.save i(vd)
x2 vd vts in2 vts ib vs ampop
XR1 GND in2 GND sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR2 in2 vd GND sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
x3 vd vts vtd GND sensor
ibias ib GND 5.53u
VSS vs GND 0
.save i(vss)
**** begin user architecture code

*cmd step stop
*PULSE ( V1 V2 TD TR TF PW PER PHASE)
.control
destroy all
save all
set color0=white
set color1=black
set temp=10
tran 10n 100u
run

plot vts out


.endc

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sym # of pins=7
** sym_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sch
.subckt sigma-delta vpwr clk out in reset_b_dff gnd vd
*.ipin in
*.iopin gnd
*.iopin clk
*.iopin out
*.iopin reset_b_dff
*.iopin vpwr
*.iopin vd
**** begin user architecture code




**** end user architecture code
XC1 in_comp gnd sky130_fd_pr__cap_mim_m3_1 W=27.196 L=27.196 MF=1 m=1
XR2 Q in_comp gnd sky130_fd_pr__res_xhigh_po_0p35 L=36 mult=1 m=1
XR1 in_comp in gnd sky130_fd_pr__res_xhigh_po_0p35 L=36 mult=1 m=1
XN1 out_comp in_comp gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XP1 out_comp in_comp vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x1 clk out_comp reset_b_dff GND GND VPWR VPWR Q out sky130_fd_sc_hd__dfrbp_1
.ends


* expanding   symbol:  /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/ampop.sym # of pins=6
** sym_path: /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/ampop.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/ampop.sch
.subckt ampop vd in1 in2 out ib vs
*.iopin vd
*.opin out
*.ipin in1
*.ipin in2
*.iopin vs
*.iopin ib
X1 vd net1 out ib vs buffer
X2 vd ib net1 in2 in1 vs ota
**** begin user architecture code


R0 in1 in1.t0 88.243
R1 in2 in2.t0 88.786
R2 vs.n0 vs.n4 362.164
R3 vs.n0 vs.n2 362.164
R4 vs.n30 vs.n25 181.834
R5 vs.n14 vs.n9 181.834
R6 vs.n18 vs.n17 108.422
R7 vs.n31 vs.n30 108.422
R8 vs.n0 vs.n6 108.422
R9 vs.n15 vs.n14 108.422
R10 vs.n34 vs.n5 5.045
R11 vs.n5 vs 0.812
R12 vs vs 0.431
R13 vs.n34 vs.n33 0.202
R14 vs vs.n34 0.182
R15 vs.n19 vs.n16 0.15
R16 vs.n32 vs.n23 0.062
R17 vs.n20 vs.n19 0.057
R18 vs.n16 vs.n7 0.055
R19 vs.n25 vs.n24 0.046
R20 vs.n9 vs.n8 0.046
R21 vs.n30 vs.n29 0.042
R22 vs.n14 vs.n13 0.042
R23 vs.n28 vs.n27 0.035
R24 vs.n12 vs.n11 0.035
R25 vs.n27 vs.n26 0.025
R26 vs.n11 vs.n10 0.025
R27 vs.n29 vs.n28 0.025
R28 vs.n13 vs.n12 0.025
R29 vs.n16 vs.n15 0.017
R30 vs.n19 vs.n18 0.017
R31 vs.n32 vs.n31 0.017
R32 vs.n4 vs.n3 0.013
R33 vs.n2 vs.n1 0.013
R34 vs.n7 vs.n0 0.007
R35 vs vs 0.005
R36 vs.n23 vs.n20 0.004
R37 vs.n33 vs.n32 0.003
R38 vs.n5 vs 0.002
R39 vs.n22 vs.n21 0.001
R40 vs.n23 vs.n22 0.001
R41 ib.n5 ib.t6 196.205
R42 ib.n6 ib.t5 196.185
R43 ib.n7 ib.t8 196.183
R44 ib.n8 ib.t7 196.181
R45 ib.n4 ib.t2 160.591
R46 ib.t2 ib.n3 160.08
R47 ib.n4 ib.t4 160.055
R48 ib.n0 ib.t9 24.837
R49 ib.n0 ib.t0 24.107
R50 ib.n1 ib.t1 17.747
R51 ib.n3 ib.t3 5.789
R52 ib.n2 ib.n1 4.041
R53 ib ib.n8 3.3
R54 ib.n5 ib.n4 1.125
R55 ib.n3 ib 0.407
R56 ib.n1 ib.n0 0.387
R57 ib.n6 ib.n5 0.175
R58 ib.n8 ib.n7 0.168
R59 ib.n7 ib.n6 0.162
R60 ib.n2 ib 0.113
R61 ib ib.n2 0.078
R62 vd.n74 vd.n73 5396.47
R63 vd.n63 vd.n62 3501.18
R64 vd.n84 vd.n83 3501.18
R65 vd.n62 vd.n59 909.81
R66 vd.n83 vd.n80 909.81
R67 vd.n65 vd.n64 722.167
R68 vd.n86 vd.n85 722.167
R69 vd.n71 vd.n70 575.623
R70 vd.n75 vd.n70 575.623
R71 vd.n74 vd.n69 569.784
R72 vd.n72 vd.n71 515.374
R73 vd.n53 vd.n52 379.482
R74 vd.n40 vd.n34 379.482
R75 vd.n61 vd.n60 373.458
R76 vd.n65 vd.n60 373.458
R77 vd.n82 vd.n81 373.458
R78 vd.n86 vd.n81 373.458
R79 vd.n69 vd.n68 326.776
R80 vd.n54 vd.n53 297.411
R81 vd.n41 vd.n40 297.411
R82 vd.n59 vd.n58 270.305
R83 vd.n80 vd.n79 270.305
R84 vd.n76 vd.n75 251.205
R85 vd.n71 vd.n68 248.846
R86 vd.n19 vd.n16 131.387
R87 vd.n4 vd.n1 131.387
R88 vd.n24 vd.n21 131.011
R89 vd.n9 vd.n6 131.011
R90 vd.n66 vd.n65 105.107
R91 vd.n87 vd.n86 105.107
R92 vd.n61 vd.n58 103.152
R93 vd.n82 vd.n79 103.152
R94 vd.n29 vd.n24 54.211
R95 vd.n14 vd.n9 54.211
R96 vd.n29 vd.n19 53.835
R97 vd.n14 vd.n4 53.835
R98 vd.n57 vd.n14 8.271
R99 vd.n57 vd.n29 7.938
R100 vd.n57 vd.n56 4.028
R101 vd.n91 vd.n90 1.897
R102 vd.n77 vd.n76 1.606
R103 vd.n67 vd.n66 1.199
R104 vd.n88 vd.n87 1.199
R105 vd.n91 vd.n57 1.058
R106 vd vd.n89 1.008
R107 vd.n78 vd.n77 0.975
R108 vd vd.n88 0.594
R109 vd.n77 vd.n68 0.389
R110 vd.n67 vd.n58 0.389
R111 vd.n88 vd.n79 0.334
R112 vd.n55 vd.n45 0.296
R113 vd.n89 vd.n78 0.273
R114 vd.n42 vd.n32 0.228
R115 vd.n56 vd.n55 0.18
R116 vd.n89 vd 0.173
R117 vd.n56 vd.n42 0.167
R118 vd.n19 vd.n18 0.161
R119 vd.n24 vd.n23 0.161
R120 vd.n4 vd.n3 0.161
R121 vd.n9 vd.n8 0.161
R122 vd.n23 vd.n22 0.139
R123 vd.n8 vd.n7 0.139
R124 vd.n18 vd.n17 0.139
R125 vd.n3 vd.n2 0.139
R126 vd.n90 vd 0.071
R127 vd.n78 vd.n67 0.054
R128 vd vd.n91 0.044
R129 vd.n90 vd 0.034
R130 vd.n42 vd.n41 0.017
R131 vd.n55 vd.n54 0.017
R132 vd.n62 vd.n61 0.015
R133 vd.n83 vd.n82 0.015
R134 vd.n16 vd.n15 0.015
R135 vd.n21 vd.n20 0.015
R136 vd.n1 vd.n0 0.015
R137 vd.n6 vd.n5 0.015
R138 vd.n52 vd.n51 0.013
R139 vd.n34 vd.n33 0.013
R140 vd.n26 vd.n25 0.013
R141 vd.n27 vd.n26 0.013
R142 vd.n11 vd.n10 0.013
R143 vd.n12 vd.n11 0.013
R144 vd.n75 vd.n74 0.004
R145 vd.n73 vd.n72 0.003
R146 vd.n63 vd.n60 0.003
R147 vd.n84 vd.n81 0.003
R148 vd.n53 vd.n50 0.003
R149 vd.n47 vd.n46 0.003
R150 vd.n36 vd.n35 0.003
R151 vd.n40 vd.n39 0.003
R152 vd.n64 vd.n63 0.003
R153 vd.n85 vd.n84 0.003
R154 vd.n50 vd.n49 0.003
R155 vd.n37 vd.n36 0.003
R156 vd.n48 vd.n47 0.003
R157 vd.n39 vd.n38 0.003
R158 vd.n73 vd.n70 0.003
R159 vd.n49 vd.n48 0.002
R160 vd.n38 vd.n37 0.002
R161 vd.n29 vd.n28 0.002
R162 vd.n28 vd.n27 0.002
R163 vd.n14 vd.n13 0.002
R164 vd.n13 vd.n12 0.002
R165 vd.n72 vd.n69 0.001
R166 vd.n64 vd.n59 0.001
R167 vd.n85 vd.n80 0.001
R168 vd.n32 vd.n31 0.001
R169 vd.n45 vd.n44 0.001
R170 vd.n44 vd.n43 0.001
R171 vd.n31 vd.n30 0.001
R172 vd.n76 vd.n69 0.001
R173 vd.n66 vd.n59 0.001
R174 vd.n87 vd.n80 0.001
R175 out.t0 out.n7 175.091
R176 out.n0 out.t2 175.044
R177 out.n2 out.n1 150.491
R178 out.n4 out.n3 150.491
R179 out.n6 out.n5 141.106
R180 out out.t0 28.743
R181 out.n5 out.t1 24.103
R182 out.n6 out.t7 24.103
R183 out.n4 out.t5 24.103
R184 out.n2 out.t3 24.102
R185 out.n0 out.t6 24.102
R186 out.n1 out.t9 24.102
R187 out.n3 out.t4 24.102
R188 out.n7 out.t8 24.102
R189 out.n7 out.n6 1.085
R190 out.n3 out.n2 0.988
R191 out.n5 out.n4 0.913
R192 out.n1 out.n0 0.863
R193 out out 0.023
R194 buffer_0/net1.n4 buffer_0/net1.t29 172.218
R195 buffer_0/net1.n5 buffer_0/net1.n4 149.523
R196 buffer_0/net1.n6 buffer_0/net1.n5 149.523
R197 buffer_0/net1.n7 buffer_0/net1.n6 149.523
R198 buffer_0/net1.n8 buffer_0/net1.n7 149.523
R199 buffer_0/net1.n9 buffer_0/net1.n8 149.523
R200 buffer_0/net1.n10 buffer_0/net1.n9 149.523
R201 buffer_0/net1.n11 buffer_0/net1.n10 149.523
R202 buffer_0/net1.n12 buffer_0/net1.n11 149.523
R203 buffer_0/net1.n13 buffer_0/net1.n12 149.523
R204 buffer_0/net1.n14 buffer_0/net1.n13 149.523
R205 buffer_0/net1.n15 buffer_0/net1.n14 149.523
R206 buffer_0/net1.n16 buffer_0/net1.n15 149.523
R207 buffer_0/net1.n17 buffer_0/net1.n16 149.523
R208 buffer_0/net1.n18 buffer_0/net1.n17 149.523
R209 buffer_0/net1.n19 buffer_0/net1.n18 149.523
R210 buffer_0/net1.n20 buffer_0/net1.n19 149.523
R211 buffer_0/net1.n21 buffer_0/net1.n20 149.523
R212 buffer_0/net1.n22 buffer_0/net1.n21 148.639
R213 buffer_0/net1.n22 buffer_0/net1.t16 24.284
R214 buffer_0/net1.n21 buffer_0/net1.t10 24.101
R215 buffer_0/net1.n20 buffer_0/net1.t27 24.101
R216 buffer_0/net1.n19 buffer_0/net1.t21 24.101
R217 buffer_0/net1.n18 buffer_0/net1.t4 24.101
R218 buffer_0/net1.n17 buffer_0/net1.t0 24.101
R219 buffer_0/net1.n16 buffer_0/net1.t22 24.101
R220 buffer_0/net1.n15 buffer_0/net1.t26 24.101
R221 buffer_0/net1.n14 buffer_0/net1.t18 24.101
R222 buffer_0/net1.n13 buffer_0/net1.t6 24.101
R223 buffer_0/net1.n12 buffer_0/net1.t23 24.101
R224 buffer_0/net1.n11 buffer_0/net1.t25 24.101
R225 buffer_0/net1.n10 buffer_0/net1.t8 24.101
R226 buffer_0/net1.n9 buffer_0/net1.t12 24.101
R227 buffer_0/net1.n8 buffer_0/net1.t28 24.101
R228 buffer_0/net1.n7 buffer_0/net1.t24 24.101
R229 buffer_0/net1.n6 buffer_0/net1.t14 24.101
R230 buffer_0/net1.n5 buffer_0/net1.t2 24.101
R231 buffer_0/net1.n4 buffer_0/net1.t20 24.101
R232 buffer_0/net1.n3 buffer_0/net1.t11 17.4
R233 buffer_0/net1.n3 buffer_0/net1.t17 17.4
R234 buffer_0/net1.n0 buffer_0/net1.t3 17.4
R235 buffer_0/net1.n0 buffer_0/net1.t15 17.4
R236 buffer_0/net1.n1 buffer_0/net1.t13 17.4
R237 buffer_0/net1.n1 buffer_0/net1.t9 17.4
R238 buffer_0/net1.n2 buffer_0/net1.t1 17.4
R239 buffer_0/net1.n2 buffer_0/net1.t5 17.4
R240 buffer_0/net1.n25 buffer_0/net1.t7 17.4
R241 buffer_0/net1.n25 buffer_0/net1.t19 17.4
R242 buffer_0/net1.n24 buffer_0/net1.n23 3.481
R243 buffer_0/net1 buffer_0/net1.n0 3.306
R244 buffer_0/net1.n27 buffer_0/net1.n26 3.218
R245 buffer_0/net1.n26 buffer_0/net1.n24 3.218
R246 buffer_0/net1.n23 buffer_0/net1.n22 1.24
R247 buffer_0/net1.n27 buffer_0/net1.n1 0.931
R248 buffer_0/net1.n24 buffer_0/net1.n2 0.931
R249 buffer_0/net1.n26 buffer_0/net1.n25 0.931
R250 buffer_0/net1 buffer_0/net1.n27 0.843
R251 buffer_0/net1.n23 buffer_0/net1.n3 0.389
C0 ota_0/m1_1300_5200# ota_0/out -0.03fF
C1 buffer_0/net2 vd 0.01fF
C2 ota_0/out vd 0.05fF
C3 buffer_0/net1.t3 vs 0.02fF
C4 buffer_0/net1.t15 vs 0.02fF
C5 buffer_0/net1.n0 vs 0.31fF $ **FLOATING
C6 buffer_0/net1.t13 vs 0.02fF
C7 buffer_0/net1.t9 vs 0.02fF
C8 buffer_0/net1.n1 vs 0.19fF $ **FLOATING
C9 buffer_0/net1.t1 vs 0.02fF
C10 buffer_0/net1.t5 vs 0.02fF
C11 buffer_0/net1.n2 vs 0.19fF $ **FLOATING
C12 buffer_0/net1.t11 vs 0.02fF
C13 buffer_0/net1.t17 vs 0.02fF
C14 buffer_0/net1.n3 vs 0.15fF $ **FLOATING
C15 buffer_0/net1.t10 vs 0.47fF
C16 buffer_0/net1.t27 vs 0.47fF
C17 buffer_0/net1.t21 vs 0.47fF
C18 buffer_0/net1.t4 vs 0.47fF
C19 buffer_0/net1.t0 vs 0.47fF
C20 buffer_0/net1.t22 vs 0.47fF
C21 buffer_0/net1.t26 vs 0.47fF
C22 buffer_0/net1.t18 vs 0.47fF
C23 buffer_0/net1.t6 vs 0.47fF
C24 buffer_0/net1.t23 vs 0.47fF
C25 buffer_0/net1.t25 vs 0.47fF
C26 buffer_0/net1.t8 vs 0.47fF
C27 buffer_0/net1.t12 vs 0.47fF
C28 buffer_0/net1.t28 vs 0.47fF
C29 buffer_0/net1.t24 vs 0.47fF
C30 buffer_0/net1.t14 vs 0.47fF
C31 buffer_0/net1.t2 vs 0.47fF
C32 buffer_0/net1.t20 vs 0.47fF
C33 buffer_0/net1.t29 vs 0.75fF
C34 buffer_0/net1.n4 vs 0.39fF $ **FLOATING
C35 buffer_0/net1.n5 vs 0.34fF $ **FLOATING
C36 buffer_0/net1.n6 vs 0.34fF $ **FLOATING
C37 buffer_0/net1.n7 vs 0.34fF $ **FLOATING
C38 buffer_0/net1.n8 vs 0.34fF $ **FLOATING
C39 buffer_0/net1.n9 vs 0.34fF $ **FLOATING
C40 buffer_0/net1.n10 vs 0.34fF $ **FLOATING
C41 buffer_0/net1.n11 vs 0.34fF $ **FLOATING
C42 buffer_0/net1.n12 vs 0.34fF $ **FLOATING
C43 buffer_0/net1.n13 vs 0.34fF $ **FLOATING
C44 buffer_0/net1.n14 vs 0.34fF $ **FLOATING
C45 buffer_0/net1.n15 vs 0.34fF $ **FLOATING
C46 buffer_0/net1.n16 vs 0.34fF $ **FLOATING
C47 buffer_0/net1.n17 vs 0.34fF $ **FLOATING
C48 buffer_0/net1.n18 vs 0.34fF $ **FLOATING
C49 buffer_0/net1.n19 vs 0.34fF $ **FLOATING
C50 buffer_0/net1.n20 vs 0.34fF $ **FLOATING
C51 buffer_0/net1.n21 vs 0.34fF $ **FLOATING
C52 buffer_0/net1.t16 vs 0.47fF
C53 buffer_0/net1.n22 vs 0.21fF $ **FLOATING
C54 buffer_0/net1.n23 vs 1.22fF $ **FLOATING
C55 buffer_0/net1.n24 vs 4.35fF $ **FLOATING
C56 buffer_0/net1.t7 vs 0.02fF
C57 buffer_0/net1.t19 vs 0.02fF
C58 buffer_0/net1.n25 vs 0.19fF $ **FLOATING
C59 buffer_0/net1.n26 vs 0.36fF $ **FLOATING
C60 buffer_0/net1.n27 vs 0.25fF $ **FLOATING
C61 out.t8 vs 0.59fF
C62 out.t1 vs 0.59fF
C63 out.t4 vs 0.59fF
C64 out.t9 vs 0.59fF
C65 out.t2 vs 0.94fF
C66 out.t6 vs 0.59fF
C67 out.n0 vs 2.69fF $ **FLOATING
C68 out.n1 vs 2.83fF $ **FLOATING
C69 out.t3 vs 0.59fF
C70 out.n2 vs 0.86fF $ **FLOATING
C71 out.n3 vs 0.86fF $ **FLOATING
C72 out.t5 vs 0.59fF
C73 out.n4 vs 0.91fF $ **FLOATING
C74 out.n5 vs 0.92fF $ **FLOATING
C75 out.t7 vs 0.59fF
C76 out.n6 vs 0.84fF $ **FLOATING
C77 out.n7 vs 0.91fF $ **FLOATING
C78 out.t0 vs 0.89fF
C79 vd.n0 vs 0.34fF $ **FLOATING
C80 vd.n1 vs 0.06fF $ **FLOATING
C81 vd.n2 vs 0.33fF $ **FLOATING
C82 vd.n3 vs 0.04fF $ **FLOATING
C83 vd.n4 vs 0.04fF $ **FLOATING
C84 vd.n5 vs 0.34fF $ **FLOATING
C85 vd.n6 vs 0.06fF $ **FLOATING
C86 vd.n7 vs 0.33fF $ **FLOATING
C87 vd.n8 vs 0.04fF $ **FLOATING
C88 vd.n9 vs 0.04fF $ **FLOATING
C89 vd.n10 vs 0.07fF $ **FLOATING
C90 vd.n11 vs 0.07fF $ **FLOATING
C91 vd.n12 vs 0.35fF $ **FLOATING
C92 vd.n13 vs 0.02fF $ **FLOATING
C93 vd.n14 vs 0.49fF $ **FLOATING
C94 vd.n15 vs 0.34fF $ **FLOATING
C95 vd.n16 vs 0.06fF $ **FLOATING
C96 vd.n17 vs 0.33fF $ **FLOATING
C97 vd.n18 vs 0.04fF $ **FLOATING
C98 vd.n19 vs 0.04fF $ **FLOATING
C99 vd.n20 vs 0.34fF $ **FLOATING
C100 vd.n21 vs 0.06fF $ **FLOATING
C101 vd.n22 vs 0.33fF $ **FLOATING
C102 vd.n23 vs 0.04fF $ **FLOATING
C103 vd.n24 vs 0.04fF $ **FLOATING
C104 vd.n25 vs 0.07fF $ **FLOATING
C105 vd.n26 vs 0.07fF $ **FLOATING
C106 vd.n27 vs 0.35fF $ **FLOATING
C107 vd.n28 vs 0.02fF $ **FLOATING
C108 vd.n29 vs 0.51fF $ **FLOATING
C109 vd.n30 vs 1.30fF $ **FLOATING
C110 vd.n31 vs 0.03fF $ **FLOATING
C111 vd.n32 vs 0.64fF $ **FLOATING
C112 vd.n33 vs 1.30fF $ **FLOATING
C113 vd.n34 vs 0.15fF $ **FLOATING
C114 vd.n35 vs 0.13fF $ **FLOATING
C115 vd.n36 vs 0.14fF $ **FLOATING
C116 vd.n37 vs 1.01fF $ **FLOATING
C117 vd.n38 vs 1.01fF $ **FLOATING
C118 vd.n39 vs 0.14fF $ **FLOATING
C119 vd.n40 vs 0.13fF $ **FLOATING
C120 vd.n41 vs 0.07fF $ **FLOATING
C121 vd.n42 vs 0.10fF $ **FLOATING
C122 vd.n43 vs 1.30fF $ **FLOATING
C123 vd.n44 vs 0.03fF $ **FLOATING
C124 vd.n45 vs 0.34fF $ **FLOATING
C125 vd.n46 vs 0.13fF $ **FLOATING
C126 vd.n47 vs 0.14fF $ **FLOATING
C127 vd.n48 vs 1.01fF $ **FLOATING
C128 vd.n49 vs 1.01fF $ **FLOATING
C129 vd.n50 vs 0.14fF $ **FLOATING
C130 vd.n51 vs 1.30fF $ **FLOATING
C131 vd.n52 vs 0.15fF $ **FLOATING
C132 vd.n53 vs 0.13fF $ **FLOATING
C133 vd.n54 vs 0.07fF $ **FLOATING
C134 vd.n55 vs 0.35fF $ **FLOATING
C135 vd.n56 vs 1.41fF $ **FLOATING
C136 vd.n57 vs 13.41fF $ **FLOATING
C137 vd.n58 vs 0.09fF $ **FLOATING
C138 vd.n59 vs 2.13fF $ **FLOATING
C139 vd.n60 vs 0.14fF $ **FLOATING
C140 vd.n61 vs 0.09fF $ **FLOATING
C141 vd.n62 vs 1.22fF $ **FLOATING
C142 vd.n63 vs 0.14fF $ **FLOATING
C143 vd.n65 vs 1.31fF $ **FLOATING
C144 vd.n66 vs 0.26fF $ **FLOATING
C145 vd.n67 vs 0.81fF $ **FLOATING
C146 vd.n68 vs 0.13fF $ **FLOATING
C147 vd.n69 vs 5.56fF $ **FLOATING
C148 vd.n70 vs 0.22fF $ **FLOATING
C149 vd.n71 vs 3.29fF $ **FLOATING
C150 vd.n73 vs 0.22fF $ **FLOATING
C151 vd.n74 vs 3.13fF $ **FLOATING
C152 vd.n75 vs 0.16fF $ **FLOATING
C153 vd.n76 vs 0.34fF $ **FLOATING
C154 vd.n77 vs 3.07fF $ **FLOATING
C155 vd.n78 vs 0.50fF $ **FLOATING
C156 vd.n79 vs 0.09fF $ **FLOATING
C157 vd.n80 vs 2.13fF $ **FLOATING
C158 vd.n81 vs 0.14fF $ **FLOATING
C159 vd.n82 vs 0.09fF $ **FLOATING
C160 vd.n83 vs 1.22fF $ **FLOATING
C161 vd.n84 vs 0.14fF $ **FLOATING
C162 vd.n86 vs 1.31fF $ **FLOATING
C163 vd.n87 vs 0.26fF $ **FLOATING
C164 vd.n88 vs 1.13fF $ **FLOATING
C165 vd.n89 vs 1.25fF $ **FLOATING
C166 vd.n90 vs 1.36fF $ **FLOATING
C167 vd.n91 vs 1.49fF $ **FLOATING
C168 ib.t1 vs 0.01fF
C169 ib.t9 vs 0.19fF
C170 ib.t0 vs 0.19fF
C171 ib.n0 vs 0.26fF $ **FLOATING
C172 ib.n1 vs 0.16fF $ **FLOATING
C173 ib.n2 vs 0.12fF $ **FLOATING
C174 ib.t8 vs 0.81fF
C175 ib.t5 vs 0.81fF
C176 ib.t6 vs 0.81fF
C177 ib.t4 vs 0.68fF
C178 ib.t3 vs 0.12fF
C179 ib.n3 vs 1.03fF $ **FLOATING
C180 ib.t2 vs 0.41fF
C181 ib.n4 vs 1.75fF $ **FLOATING
C182 ib.n5 vs 0.99fF $ **FLOATING
C183 ib.n6 vs 0.51fF $ **FLOATING
C184 ib.n7 vs 0.52fF $ **FLOATING
C185 ib.t7 vs 0.81fF
C186 ib.n8 vs 1.32fF $ **FLOATING
C187 buffer_0/net4 vs 1.11fF
C188 out vs 13.18fF
C189 buffer_0/net3 vs 2.90fF
C190 vd vs 38.03fF
C191 buffer_0/net1 vs 14.70fF
C192 buffer_0/net2 vs 3.06fF
C193 ota_0/out vs 11.16fF
C194 ota_0/m1_n20_5200# vs 2.40fF
C195 ota_0/m1_420_6300# vs 4.72fF
C196 ota_0/m1_1300_5200# vs 14.02fF


**** end user architecture code
.ends


* expanding   symbol:  /home/hugodg/projects-sky130/temp-sensor/sensor/xschem/sensor.sym # of pins=4
** sym_path: /home/hugodg/projects-sky130/temp-sensor/sensor/xschem/sensor.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/sensor/xschem/sensor.sch
.subckt sensor vd vts vtd gnd
*.iopin vd
*.opin vts
*.opin vtd
*.iopin gnd
XP1 a a vd vd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP2 c a d d sky130_fd_pr__pfet_01v8 L=1 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP3 d vtd vd vd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP4 vts vtd vd vd sky130_fd_pr__pfet_01v8 L=5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP5 b vtd c c sky130_fd_pr__pfet_01v8 L=1 W=8 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP6 vtd vtd vts vts sky130_fd_pr__pfet_01v8 L=1 W=16 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XN1 a b gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XN2 b b gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XN3 vtd b gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
**** begin user architecture code


R0 vd.n23 vd.n22 222.87
R1 vd.n10 vd.n9 222.87
R2 vd.n24 vd.n23 149.458
R3 vd.n11 vd.n10 149.458
R4 vd.n26 vd.n12 0.85
R5 vd.n26 vd.n25 0.375
R6 vd.n25 vd.n15 0.37
R7 vd.n12 vd.n2 0.37
R8 vd vd.n26 0.112
R9 vd.n25 vd.n24 0.017
R10 vd.n12 vd.n11 0.017
R11 vd.n22 vd.n21 0.015
R12 vd.n9 vd.n8 0.015
R13 vd.n23 vd.n20 0.008
R14 vd.n17 vd.n16 0.008
R15 vd.n10 vd.n7 0.008
R16 vd.n4 vd.n3 0.008
R17 vd.n20 vd.n19 0.006
R18 vd.n7 vd.n6 0.006
R19 vd.n18 vd.n17 0.006
R20 vd.n5 vd.n4 0.006
R21 vd.n19 vd.n18 0.004
R22 vd.n6 vd.n5 0.004
R23 vd.n15 vd.n14 0.001
R24 vd.n2 vd.n1 0.001
R25 vd.n14 vd.n13 0.001
R26 vd.n1 vd.n0 0.001
R27 vtd.n19 vtd.t21 64.503
R28 vtd.n1 vtd.t20 63.858
R29 vtd.n11 vtd.t0 63.734
R30 vtd.n17 vtd.t18 63.628
R31 vtd.n16 vtd.t17 63.628
R32 vtd.n15 vtd.t2 63.628
R33 vtd.n13 vtd.t4 63.628
R34 vtd.n12 vtd.t6 63.628
R35 vtd.n8 vtd.t8 63.628
R36 vtd.n4 vtd.t12 63.628
R37 vtd.n5 vtd.t14 63.628
R38 vtd.n1 vtd.t19 63.628
R39 vtd.n2 vtd.t10 63.628
R40 vtd.n10 vtd.t1 14.282
R41 vtd.n10 vtd.t7 14.282
R42 vtd.n9 vtd.t5 14.282
R43 vtd.n9 vtd.t3 14.282
R44 vtd.n6 vtd.t9 14.282
R45 vtd.n6 vtd.t15 14.282
R46 vtd.n0 vtd.t13 14.282
R47 vtd.n0 vtd.t11 14.282
R48 vtd.n19 vtd.t16 12.724
R49 vtd.n2 vtd.n1 0.787
R50 vtd.n16 vtd.n15 0.769
R51 vtd vtd.n20 0.568
R52 vtd.n18 vtd.n17 0.478
R53 vtd.n20 vtd.n18 0.244
R54 vtd.n17 vtd.n16 0.23
R55 vtd.n20 vtd.n19 0.16
R56 vtd.n8 vtd.n7 0.105
R57 vtd.n15 vtd.n14 0.1
R58 vtd.n3 vtd.n2 0.1
R59 vtd.n13 vtd.n12 0.089
R60 vtd.n5 vtd.n4 0.089
R61 vtd.n18 vtd.n8 0.08
R62 vtd.n11 vtd.n10 0.061
R63 vtd.n7 vtd.n6 0.061
R64 vtd.n14 vtd.n9 0.057
R65 vtd.n3 vtd.n0 0.057
R66 vtd.n12 vtd.n11 0.045
R67 vtd.n7 vtd.n5 0.045
R68 vtd.n14 vtd.n13 0.044
R69 vtd.n4 vtd.n3 0.044
R70 vts.n6 vts.n5 151.046
R71 vts.n8 vts.n7 149.458
R72 vts vts.n9 2.772
R73 vts.n9 vts.n6 1.514
R74 vts.n9 vts.n8 0.017
R75 vts.n5 vts.n4 0.008
R76 vts.n1 vts.n0 0.004
R77 vts.n2 vts.n1 0.004
R78 vts.n3 vts.n2 0.001
R79 vts.n6 vts.n3 0.001
R80 b.n1 b.t7 17.619
R81 b.n7 b.t4 18.027
R82 b.n0 b.t3 17.404
R83 b.n2 b.t2 17.404
R84 b.n2 b.t6 18.003
R85 b.n11 b.t0 17.404
R86 b.n9 b.t5 17.404
R87 b.n7 b.t1 17.404
R88 b.n19 b.n12 6.22
R89 b.n16 b.n15 4.5
R90 b.n16 b.n14 4.5
R91 b.n4 b.n1 3.868
R92 b.n4 b.n3 3.839
R93 b.n17 b.n16 2.625
R94 b.n6 b.n5 1.507
R95 b b.n19 0.928
R96 b.n6 b.n4 0.708
R97 b.n19 b.n6 0.708
R98 b.n18 b.n17 0.708
R99 b.n19 b.n18 0.666
R100 b.n9 b.n8 0.45
R101 b.n11 b.n10 0.448
R102 b.n1 b.n0 0.356
R103 b.n12 b.n11 0.17
R104 b.n10 b.n9 0.168
R105 b.n3 b.n2 0.16
R106 b.n8 b.n7 0.159
R107 b.n14 b.n13 0.113
R108 gnd.n0 gnd.n5 732.611
R109 gnd.n0 gnd.n3 732.611
R110 gnd.n34 gnd.n33 732.611
R111 gnd.n34 gnd.n10 732.611
R112 gnd.n44 gnd.n43 732.611
R113 gnd.n44 gnd.n40 732.611
R114 gnd.n10 gnd.n8 659.199
R115 gnd.n40 gnd.n38 659.199
R116 gnd.n33 gnd.n31 653.176
R117 gnd.n43 gnd.n41 649.411
R118 gnd.n30 gnd.n16 31.079
R119 gnd.n8 gnd.n7 30.494
R120 gnd.n16 gnd.n11 19.019
R121 gnd.n23 gnd.n22 9.3
R122 gnd.n16 gnd.n15 9.3
R123 gnd.n20 gnd.n19 9.3
R124 gnd.n38 gnd.n35 7.529
R125 gnd.n49 gnd.n48 7.152
R126 gnd.n31 gnd.n30 6.023
R127 gnd.n6 gnd.n57 2.258
R128 gnd.n0 gnd.n21 1.876
R129 gnd.n66 gnd.n65 0.186
R130 gnd.n64 gnd.n63 0.18
R131 gnd.n59 gnd.n58 0.107
R132 gnd.n27 gnd.n26 0.102
R133 gnd.n24 gnd.n20 0.077
R134 gnd.n15 gnd.n14 0.072
R135 gnd gnd.n1 0.07
R136 gnd.n66 gnd.n62 0.069
R137 gnd.n0 gnd.n23 0.067
R138 gnd.n28 gnd.n27 0.066
R139 gnd.n37 gnd.n36 0.062
R140 gnd.n25 gnd.n18 0.056
R141 gnd.n1 gnd.n70 0.055
R142 gnd.n60 gnd.n56 0.052
R143 gnd.n61 gnd.n60 0.046
R144 gnd.n1 gnd.n67 0.046
R145 gnd.n59 gnd.n6 0.046
R146 gnd.n24 gnd.n0 0.046
R147 gnd.n1 gnd.n34 0.046
R148 gnd.n6 gnd.n44 0.046
R149 gnd.n1 gnd.n69 0.045
R150 gnd.n29 gnd.n17 0.039
R151 gnd.n29 gnd.n28 0.039
R152 gnd.n67 gnd.n45 0.034
R153 gnd.n61 gnd.n51 0.034
R154 gnd.n15 gnd.n12 0.031
R155 gnd.n55 gnd.n53 0.03
R156 gnd.n30 gnd.n29 0.03
R157 gnd.n51 gnd.n50 0.025
R158 gnd.n14 gnd.n13 0.023
R159 gnd.n60 gnd.n59 0.019
R160 gnd.n50 gnd.n47 0.018
R161 gnd.n38 gnd.n37 0.017
R162 gnd.n50 gnd.n49 0.017
R163 gnd.n66 gnd.n64 0.012
R164 gnd.n53 gnd.n52 0.011
R165 gnd.n56 gnd.n55 0.01
R166 gnd.n26 gnd.n25 0.009
R167 gnd.n25 gnd.n24 0.006
R168 gnd.n69 gnd.n68 0.005
R169 gnd.n5 gnd.n4 0.004
R170 gnd.n3 gnd.n2 0.004
R171 gnd.n33 gnd.n32 0.004
R172 gnd.n10 gnd.n9 0.004
R173 gnd.n43 gnd.n42 0.004
R174 gnd.n40 gnd.n39 0.004
R175 gnd.n55 gnd.n54 0.002
R176 gnd.n67 gnd.n66 0.001
R177 gnd.n62 gnd.n61 0.001
R178 gnd.n62 gnd.n46 0.001
C0 vts vtd 7.80fF
C1 b c 2.09fF
C2 vd vtd 2.64fF
C3 vtd c 3.54fF
C4 vtd b 5.31fF
C5 a d 4.24fF
C6 a vts 0.90fF
C7 a vd 0.99fF
C8 a c 1.42fF
C9 a b 4.95fF
C10 d vts 0.21fF
C11 d vd 1.91fF
C12 a vtd 1.18fF
C13 d c 1.52fF
C14 d b 0.38fF
C15 d vtd 0.54fF
C16 vd vts 0.43fF
C17 vts c 1.96fF
C18 vts b 4.21fF
C19 vd c 0.64fF
C20 vd b 0.24fF
C21 b.t7 gnd 0.15fF
C22 b.t3 gnd 0.10fF
C23 b.n0 gnd 2.66fF $ **FLOATING
C24 b.n1 gnd 7.23fF $ **FLOATING
C25 b.t6 gnd 0.18fF
C26 b.t2 gnd 0.10fF
C27 b.n2 gnd 3.85fF $ **FLOATING
C28 b.n3 gnd 3.44fF $ **FLOATING
C29 b.n4 gnd 14.60fF $ **FLOATING
C30 b.n5 gnd 4.96fF $ **FLOATING
C31 b.n6 gnd 2.62fF $ **FLOATING
C32 b.t4 gnd 0.17fF
C33 b.t1 gnd 0.10fF
C34 b.n7 gnd 3.24fF $ **FLOATING
C35 b.n8 gnd 2.43fF $ **FLOATING
C36 b.t5 gnd 0.10fF
C37 b.n9 gnd 1.17fF $ **FLOATING
C38 b.n10 gnd 2.45fF $ **FLOATING
C39 b.t0 gnd 0.10fF
C40 b.n11 gnd 1.19fF $ **FLOATING
C41 b.n12 gnd 2.60fF $ **FLOATING
C42 b.n13 gnd 0.26fF $ **FLOATING
C43 b.n14 gnd 0.19fF $ **FLOATING
C44 b.n15 gnd 0.08fF $ **FLOATING
C45 b.n16 gnd 4.36fF $ **FLOATING
C46 b.n17 gnd 7.09fF $ **FLOATING
C47 b.n18 gnd 5.66fF $ **FLOATING
C48 b.n19 gnd 7.78fF $ **FLOATING
C49 vts.n0 gnd 0.19fF $ **FLOATING
C50 vts.n1 gnd 0.19fF $ **FLOATING
C51 vts.n3 gnd 3.30fF $ **FLOATING
C52 vts.n4 gnd 1.95fF $ **FLOATING
C53 vts.n5 gnd 0.14fF $ **FLOATING
C54 vts.n6 gnd 0.33fF $ **FLOATING
C55 vts.n7 gnd 2.08fF $ **FLOATING
C56 vts.n8 gnd 0.10fF $ **FLOATING
C57 vts.n9 gnd 8.26fF $ **FLOATING
C58 vtd.t8 gnd 0.47fF
C59 vtd.t14 gnd 0.47fF
C60 vtd.t12 gnd 0.47fF
C61 vtd.t13 gnd 0.03fF
C62 vtd.t11 gnd 0.03fF
C63 vtd.n0 gnd 0.13fF $ **FLOATING
C64 vtd.t10 gnd 0.47fF
C65 vtd.t19 gnd 0.47fF
C66 vtd.t20 gnd 0.47fF
C67 vtd.n1 gnd 0.89fF $ **FLOATING
C68 vtd.n2 gnd 0.51fF $ **FLOATING
C69 vtd.n3 gnd 0.18fF $ **FLOATING
C70 vtd.n4 gnd 0.51fF $ **FLOATING
C71 vtd.n5 gnd 0.51fF $ **FLOATING
C72 vtd.t9 gnd 0.03fF
C73 vtd.t15 gnd 0.03fF
C74 vtd.n6 gnd 0.13fF $ **FLOATING
C75 vtd.n7 gnd 0.18fF $ **FLOATING
C76 vtd.n8 gnd 0.25fF $ **FLOATING
C77 vtd.t5 gnd 0.03fF
C78 vtd.t3 gnd 0.03fF
C79 vtd.n9 gnd 0.13fF $ **FLOATING
C80 vtd.t0 gnd 0.47fF
C81 vtd.t1 gnd 0.03fF
C82 vtd.t7 gnd 0.03fF
C83 vtd.n10 gnd 0.13fF $ **FLOATING
C84 vtd.n11 gnd 0.46fF $ **FLOATING
C85 vtd.t6 gnd 0.47fF
C86 vtd.n12 gnd 0.51fF $ **FLOATING
C87 vtd.t4 gnd 0.47fF
C88 vtd.n13 gnd 0.51fF $ **FLOATING
C89 vtd.n14 gnd 0.18fF $ **FLOATING
C90 vtd.t2 gnd 0.47fF
C91 vtd.n15 gnd 0.50fF $ **FLOATING
C92 vtd.t17 gnd 0.47fF
C93 vtd.n16 gnd 0.55fF $ **FLOATING
C94 vtd.t18 gnd 0.47fF
C95 vtd.n17 gnd 0.44fF $ **FLOATING
C96 vtd.n18 gnd 0.54fF $ **FLOATING
C97 vtd.t16 gnd 2.35fF
C98 vtd.t21 gnd 0.48fF
C99 vtd.n19 gnd 2.32fF $ **FLOATING
C100 vtd.n20 gnd 7.12fF $ **FLOATING
C101 vd.n0 gnd 0.62fF $ **FLOATING
C102 vd.n1 gnd 0.03fF $ **FLOATING
C103 vd.n2 gnd 0.09fF $ **FLOATING
C104 vd.n3 gnd 0.07fF $ **FLOATING
C105 vd.n4 gnd 0.08fF $ **FLOATING
C106 vd.n5 gnd 0.42fF $ **FLOATING
C107 vd.n6 gnd 0.42fF $ **FLOATING
C108 vd.n7 gnd 0.08fF $ **FLOATING
C109 vd.n8 gnd 0.62fF $ **FLOATING
C110 vd.n9 gnd 0.08fF $ **FLOATING
C111 vd.n10 gnd 0.07fF $ **FLOATING
C112 vd.n11 gnd 0.04fF $ **FLOATING
C113 vd.n12 gnd 0.98fF $ **FLOATING
C114 vd.n13 gnd 0.62fF $ **FLOATING
C115 vd.n14 gnd 0.03fF $ **FLOATING
C116 vd.n15 gnd 0.09fF $ **FLOATING
C117 vd.n16 gnd 0.07fF $ **FLOATING
C118 vd.n17 gnd 0.08fF $ **FLOATING
C119 vd.n18 gnd 0.42fF $ **FLOATING
C120 vd.n19 gnd 0.42fF $ **FLOATING
C121 vd.n20 gnd 0.08fF $ **FLOATING
C122 vd.n21 gnd 0.62fF $ **FLOATING
C123 vd.n22 gnd 0.08fF $ **FLOATING
C124 vd.n23 gnd 0.07fF $ **FLOATING
C125 vd.n24 gnd 0.04fF $ **FLOATING
C126 vd.n25 gnd 14.58fF $ **FLOATING
C127 vd.n26 gnd 3.50fF $ **FLOATING
C128 d gnd 9.68fF
C129 a gnd 10.08fF
C130 c gnd -15.39fF
C131 b gnd 131.16fF
C132 vtd gnd -35.85fF
C133 vts gnd 18.71fF
C134 vd gnd 13.44fF


**** end user architecture code
.ends


* expanding   symbol:  /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/buffer.sym # of pins=5
** sym_path: /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/buffer.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/buffer.sch
.subckt buffer vd in out ib gnd
*.iopin vd
*.iopin ib
*.iopin out
*.iopin in
*.iopin gnd
XM3 net2 net2 vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 out net4 gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 in net4 gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 net3 vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 ib gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out net3 vd vd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out net1 gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net1 net2 vd vd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 net1 gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 ib ib gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/ota.sym # of pins=6
** sym_path: /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/ota.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/amp-op/xschem/ota.sch
.subckt ota vd ib out in2 in1 vs
*.iopin vd
*.iopin vs
*.iopin ib
*.ipin in1
*.ipin in2
*.opin out
XCC out d sky130_fd_pr__cap_mim_m3_1 W=21 L=21 MF=1 m=1
XM5 ib ib vd vd sky130_fd_pr__pfet_01v8 L=1 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 b ib vd vd sky130_fd_pr__pfet_01v8 L=1 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 out ib vd vd sky130_fd_pr__pfet_01v8 L=1 W=30 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 c in1 b b sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 d in2 b b sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 c c vs vs sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 d c vs vs sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out d vs vs sky130_fd_pr__nfet_01v8 L=1 W=9 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
