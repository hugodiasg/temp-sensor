magic
tech sky130A
magscale 1 2
timestamp 1675640756
<< psubdiff >>
rect 4776 4200 4800 4700
rect 5700 4200 5724 4700
<< psubdiffcont >>
rect 4800 4200 5700 4700
<< locali >>
rect 4784 4200 4800 4700
rect 5700 4200 5716 4700
<< viali >>
rect 4800 4200 5700 4700
<< metal1 >>
rect -28700 7200 -21200 7300
rect -28700 5700 -22600 7200
rect -21400 5700 -21200 7200
rect -28700 5600 -21200 5700
rect -28700 5500 -21300 5600
rect 3500 4700 6400 4800
rect 3500 4200 3600 4700
rect 4600 4200 4800 4700
rect 5700 4200 6400 4700
rect 3500 4100 6400 4200
rect 2000 -11700 6500 -11600
rect 1900 -11800 6500 -11700
rect 1900 -13300 2100 -11800
rect 3300 -13300 6500 -11800
rect 1900 -13400 6500 -13300
<< via1 >>
rect -22600 5700 -21400 7200
rect 3600 4200 4600 4700
rect 2100 -13300 3300 -11800
<< metal2 >>
rect -22700 7200 -21200 7300
rect -22700 5700 -22600 7200
rect -21400 5700 -21200 7200
rect -22700 5600 -21200 5700
rect 3500 4700 4700 4800
rect 3500 4200 3600 4700
rect 4600 4200 4700 4700
rect 3500 4100 4700 4200
rect 1900 -11800 3400 -11700
rect 1900 -13300 2100 -11800
rect 3300 -13300 3400 -11800
rect 1900 -13400 3400 -13300
<< via2 >>
rect -22600 5700 -21400 7200
rect 3600 4200 4600 4700
rect 2100 -13300 3300 -11800
<< metal3 >>
rect -22700 7200 -21200 7300
rect -22700 5700 -22600 7200
rect -21400 5700 -21200 7200
rect -22700 5600 -21200 5700
rect 3500 4700 4700 4800
rect 3500 4200 3600 4700
rect 4600 4200 4700 4700
rect 3500 4100 4700 4200
rect 1900 -11800 3400 -11700
rect 1900 -13300 2100 -11800
rect 3300 -13300 3400 -11800
rect 1900 -13400 3400 -13300
<< via3 >>
rect -22600 5700 -21400 7200
rect 3600 4200 4600 4700
rect 2100 -13300 3300 -11800
<< metal4 >>
rect -22744 7222 -21184 7328
rect -22744 5588 -22604 7222
rect -21358 5588 -21184 7222
rect -22744 4582 -21184 5588
rect -16047 5435 -15685 5485
rect -16286 5402 -15685 5435
rect -19058 4646 -15652 5402
rect -13348 4646 -10468 5978
rect -8722 4646 -5546 5798
rect -4130 4646 -198 6488
rect 938 5100 4938 6818
rect 938 4700 4800 5100
rect 938 4646 3600 4700
rect -22744 2810 -21172 4582
rect -19058 4300 3600 4646
rect -16286 4284 3600 4300
rect -11560 3406 -6680 4284
rect -5656 3176 -1204 4284
rect 50 4200 3600 4284
rect 4600 4284 4800 4700
rect 4600 4200 4798 4284
rect 50 3044 4798 4200
rect 1900 -11688 3444 -11600
rect 1900 -13322 2058 -11688
rect 3304 -13322 3444 -11688
rect 1900 -13428 3444 -13322
<< via4 >>
rect -22604 7200 -21358 7222
rect -22604 5700 -22600 7200
rect -22600 5700 -21400 7200
rect -21400 5700 -21358 7200
rect -22604 5588 -21358 5700
rect 2058 -11800 3304 -11688
rect 2058 -13300 2100 -11800
rect 2100 -13300 3300 -11800
rect 3300 -13300 3304 -11800
rect 2058 -13322 3304 -13300
<< metal5 >>
rect -17250 27020 3100 28804
rect -17250 25444 -15466 27020
rect -13294 25184 -11510 27020
rect -7924 25054 -6140 27020
rect -3142 25184 -1358 27020
rect 1316 25672 3100 27020
rect -22734 7282 -21174 7328
rect -22734 7222 -16936 7282
rect -22734 5588 -22604 7222
rect -21358 5588 -16936 7222
rect -22734 5498 -16936 5588
rect -22734 5476 -21174 5498
rect -10079 -11618 -8509 -10029
rect -4223 -11618 -2653 -10159
rect 1635 -11600 3205 -9277
rect 1635 -11618 3434 -11600
rect -14431 -11688 3434 -11618
rect -14431 -13188 2058 -11688
rect 1900 -13322 2058 -13188
rect 3304 -13322 3434 -11688
rect 1900 -13428 3434 -13322
use 1  1_0
timestamp 1675570359
transform -1 0 30546 0 -1 46012
box 43200 41630 59200 59200
use sky130_fd_pr__cap_mim_m3_2_MH6WNN  XC0
timestamp 1675569099
transform 1 0 -3067 0 1 -3500
box -8407 -7560 8429 7560
use sky130_fd_pr__cap_mim_m3_2_C96Y74  XC1
timestamp 1675569099
transform 1 0 -6887 0 1 15834
box -12345 -10800 12367 10800
<< labels >>
flabel metal1 5800 4100 6400 4800 0 FreeSans 8000 0 0 0 gnd
port 2 nsew
flabel metal1 -28700 5500 -27600 7300 0 FreeSans 8000 0 0 0 out
port 4 nsew
flabel metal1 5400 -13400 6500 -11600 0 FreeSans 8000 0 0 0 in
port 6 nsew
<< end >>
