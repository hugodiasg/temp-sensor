magic
tech sky130A
timestamp 1646185352
<< metal4 >>
rect 25805 26581 30394 26600
rect 25805 25823 25823 26581
rect 26581 25823 30394 26581
rect 25805 25805 30394 25823
<< via4 >>
rect 25823 25823 26581 26581
<< metal5 >>
rect 21600 28805 29600 29600
rect 21600 27805 28600 28600
rect 21600 22394 22394 27805
rect 22599 26805 27600 27600
rect 22599 23394 23394 26805
rect 23599 26581 26600 26600
rect 23599 25823 25823 26581
rect 26581 25823 26600 26581
rect 23599 25805 26600 25823
rect 23599 24394 24394 25805
rect 26805 24394 27600 26805
rect 23599 23599 27600 24394
rect 27805 23394 28600 27805
rect 22599 22599 28600 23394
rect 28805 22394 29600 28805
rect 21600 21600 29600 22394
<< end >>
