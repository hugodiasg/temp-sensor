magic
tech sky130A
magscale 1 2
timestamp 1646425662
<< metal4 >>
rect -2609 7649 2609 7690
rect -2609 2671 2353 7649
rect 2589 2671 2609 7649
rect -2609 2630 2609 2671
rect -2609 2489 2609 2530
rect -2609 -2489 2353 2489
rect 2589 -2489 2609 2489
rect -2609 -2530 2609 -2489
rect -2609 -2671 2609 -2630
rect -2609 -7649 2353 -2671
rect 2589 -7649 2609 -2671
rect -2609 -7690 2609 -7649
<< via4 >>
rect 2353 2671 2589 7649
rect 2353 -2489 2589 2489
rect 2353 -7649 2589 -2671
<< mimcap2 >>
rect -2509 7550 2351 7590
rect -2509 2770 -1991 7550
rect 1833 2770 2351 7550
rect -2509 2730 2351 2770
rect -2509 2390 2351 2430
rect -2509 -2390 -1991 2390
rect 1833 -2390 2351 2390
rect -2509 -2430 2351 -2390
rect -2509 -2770 2351 -2730
rect -2509 -7550 -1991 -2770
rect 1833 -7550 2351 -2770
rect -2509 -7590 2351 -7550
<< mimcap2contact >>
rect -1991 2770 1833 7550
rect -1991 -2390 1833 2390
rect -1991 -7550 1833 -2770
<< metal5 >>
rect -239 7574 81 7740
rect 2311 7649 2631 7740
rect -2015 7550 1857 7574
rect -2015 2770 -1991 7550
rect 1833 2770 1857 7550
rect -2015 2746 1857 2770
rect -239 2414 81 2746
rect 2311 2671 2353 7649
rect 2589 2671 2631 7649
rect 2311 2489 2631 2671
rect -2015 2390 1857 2414
rect -2015 -2390 -1991 2390
rect 1833 -2390 1857 2390
rect -2015 -2414 1857 -2390
rect -239 -2746 81 -2414
rect 2311 -2489 2353 2489
rect 2589 -2489 2631 2489
rect 2311 -2671 2631 -2489
rect -2015 -2770 1857 -2746
rect -2015 -7550 -1991 -2770
rect 1833 -7550 1857 -2770
rect -2015 -7574 1857 -7550
rect -239 -7740 81 -7574
rect 2311 -7649 2353 -2671
rect 2589 -7649 2631 -2671
rect 2311 -7740 2631 -7649
<< properties >>
string FIXED_BBOX -2609 2630 2451 7690
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.3 l 24.3 val 1.199k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
