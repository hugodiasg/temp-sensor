** sch_path: /foss/designs/temp-sensor/buffer/xschem/buffer.sch
.subckt buffer vd ib out in gnd
*.PININFO vd:B ib:B out:B in:B gnd:B
XM3 a a vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM1 a out c gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 m=1
XM2 b in c gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 m=1
XM4 b b vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM5 c ib gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM6 out b vd vd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=10 m=1
XM7 out d gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 m=1
XM8 d a vd vd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=10 m=1
XM9 d d gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 m=1
XM10 ib ib gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XCc out d sky130_fd_pr__cap_mim_m3_2 W=30 L=15 m=1
XM11 vd vd vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM12 vd vd vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM13 a a a gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM14 a a a gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM15 ib ib ib gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM16 d d d gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends
.end
