magic
tech sky130A
magscale 1 2
timestamp 1646014094
<< metal4 >>
rect -2681 10517 2681 10558
rect -2681 5395 2425 10517
rect 2661 5395 2681 10517
rect -2681 5354 2681 5395
rect -2681 5213 2681 5254
rect -2681 91 2425 5213
rect 2661 91 2681 5213
rect -2681 50 2681 91
rect -2681 -91 2681 -50
rect -2681 -5213 2425 -91
rect 2661 -5213 2681 -91
rect -2681 -5254 2681 -5213
rect -2681 -5395 2681 -5354
rect -2681 -10517 2425 -5395
rect 2661 -10517 2681 -5395
rect -2681 -10558 2681 -10517
<< via4 >>
rect 2425 5395 2661 10517
rect 2425 91 2661 5213
rect 2425 -5213 2661 -91
rect 2425 -10517 2661 -5395
<< mimcap2 >>
rect -2581 10418 2423 10458
rect -2581 5494 -2049 10418
rect 1891 5494 2423 10418
rect -2581 5454 2423 5494
rect -2581 5114 2423 5154
rect -2581 190 -2049 5114
rect 1891 190 2423 5114
rect -2581 150 2423 190
rect -2581 -190 2423 -150
rect -2581 -5114 -2049 -190
rect 1891 -5114 2423 -190
rect -2581 -5154 2423 -5114
rect -2581 -5494 2423 -5454
rect -2581 -10418 -2049 -5494
rect 1891 -10418 2423 -5494
rect -2581 -10458 2423 -10418
<< mimcap2contact >>
rect -2049 5494 1891 10418
rect -2049 190 1891 5114
rect -2049 -5114 1891 -190
rect -2049 -10418 1891 -5494
<< metal5 >>
rect -239 10442 81 10608
rect 2383 10517 2703 10608
rect -2073 10418 1915 10442
rect -2073 5494 -2049 10418
rect 1891 5494 1915 10418
rect -2073 5470 1915 5494
rect -239 5138 81 5470
rect 2383 5395 2425 10517
rect 2661 5395 2703 10517
rect 2383 5213 2703 5395
rect -2073 5114 1915 5138
rect -2073 190 -2049 5114
rect 1891 190 1915 5114
rect -2073 166 1915 190
rect -239 -166 81 166
rect 2383 91 2425 5213
rect 2661 91 2703 5213
rect 2383 -91 2703 91
rect -2073 -190 1915 -166
rect -2073 -5114 -2049 -190
rect 1891 -5114 1915 -190
rect -2073 -5138 1915 -5114
rect -239 -5470 81 -5138
rect 2383 -5213 2425 -91
rect 2661 -5213 2703 -91
rect 2383 -5395 2703 -5213
rect -2073 -5494 1915 -5470
rect -2073 -10418 -2049 -5494
rect 1891 -10418 1915 -5494
rect -2073 -10442 1915 -10418
rect -239 -10608 81 -10442
rect 2383 -10517 2425 -5395
rect 2661 -10517 2703 -5395
rect 2383 -10608 2703 -10517
<< properties >>
string FIXED_BBOX -2681 5354 2523 10558
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.019 l 25.019 val 1.27k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
