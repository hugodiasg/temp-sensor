magic
tech sky130A
magscale 1 2
timestamp 1700108998
<< metal4 >>
rect -2789 7759 2789 7800
rect -2789 2801 2533 7759
rect 2769 2801 2789 7759
rect -2789 2760 2789 2801
rect -2789 2479 2789 2520
rect -2789 -2479 2533 2479
rect 2769 -2479 2789 2479
rect -2789 -2520 2789 -2479
rect -2789 -2801 2789 -2760
rect -2789 -7759 2533 -2801
rect 2769 -7759 2789 -2801
rect -2789 -7800 2789 -7759
<< via4 >>
rect 2533 2801 2769 7759
rect 2533 -2479 2769 2479
rect 2533 -7759 2769 -2801
<< mimcap2 >>
rect -2709 7680 2171 7720
rect -2709 2880 -2669 7680
rect 2131 2880 2171 7680
rect -2709 2840 2171 2880
rect -2709 2400 2171 2440
rect -2709 -2400 -2669 2400
rect 2131 -2400 2171 2400
rect -2709 -2440 2171 -2400
rect -2709 -2880 2171 -2840
rect -2709 -7680 -2669 -2880
rect 2131 -7680 2171 -2880
rect -2709 -7720 2171 -7680
<< mimcap2contact >>
rect -2669 2880 2131 7680
rect -2669 -2400 2131 2400
rect -2669 -7680 2131 -2880
<< metal5 >>
rect -429 7704 -109 7920
rect 2491 7759 2811 7920
rect -2693 7680 2155 7704
rect -2693 2880 -2669 7680
rect 2131 2880 2155 7680
rect -2693 2856 2155 2880
rect -429 2424 -109 2856
rect 2491 2801 2533 7759
rect 2769 2801 2811 7759
rect 2491 2479 2811 2801
rect -2693 2400 2155 2424
rect -2693 -2400 -2669 2400
rect 2131 -2400 2155 2400
rect -2693 -2424 2155 -2400
rect -429 -2856 -109 -2424
rect 2491 -2479 2533 2479
rect 2769 -2479 2811 2479
rect 2491 -2801 2811 -2479
rect -2693 -2880 2155 -2856
rect -2693 -7680 -2669 -2880
rect 2131 -7680 2155 -2880
rect -2693 -7704 2155 -7680
rect -429 -7920 -109 -7704
rect 2491 -7759 2533 -2801
rect 2769 -7759 2811 -2801
rect 2491 -7920 2811 -7759
<< properties >>
string FIXED_BBOX -2789 2760 2251 7800
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.4 l 24.4 val 1.209k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
