* NGSPICE file created from buffer.ext - technology: sky130A

.subckt buffer vd ib out in gnd
X0 b.t12 b.t11 vd.t18 vd.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 vd.t25 vd.t22 vd.t24 vd.t23 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X2 c out a gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X3 out.t7 d.t12 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a a a vd.t41 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=1.16 ps=10.3 w=1 l=1
X5 d.t11 a vd.t40 vd.t39 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X6 d.t5 d.t4 d.t5 vd.t42 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0 w=15 l=1
X7 vd.t21 vd.t19 vd.t21 vd.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X8 a a vd.t38 vd.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X9 gnd.t24 d.t13 out.t8 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 vd.t16 b.t16 out.t6 vd.t15 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X11 out.t4 out.t2 out.t3 vd.t0 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0 w=15 l=1
X12 d.t9 d.t8 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a a vd.t36 vd.t35 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 b.t6 b.t4 b.t5 vd.t14 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X15 a a a gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0.96 ps=7.28 w=1.5 l=0.15
X16 gnd.t20 gnd.t17 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=1
X17 vd.t34 a a vd.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 vd.t32 a a vd.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 a a vd.t30 vd.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 b.t3 b.t2 b.t3 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0 ps=0 w=1.5 l=0.15
X21 gnd.t1 ib.t3 ib.t4 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 c ib.t5 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 ib.t2 ib.t0 ib.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X24 out.t5 b.t17 vd.t13 vd.t12 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X25 b.t10 b.t9 vd vd.t9 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 vd b.t7 b.t8 vd.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 gnd.t22 d.t6 d.t7 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 out.t1 out.t0 out.t1 vd.t26 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0 w=15 l=1
X29 vd.t5 b.t13 b.t14 vd.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X30 b.t15 in.t0 c gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X31 c c c gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=1.08 ps=8.82 w=1 l=1
X32 vd.t28 a d.t10 vd.t27 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X33 d.t3 d.t1 d.t2 vd.t1 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0 w=15 l=1
X34 out d.t0 sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X35 vd.t3 b.t0 b.t1 vd.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 gnd.t16 gnd.t14 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=1
R0 b.n11 b.t17 377.466
R1 b.n11 b.t16 376.93
R2 b.n18 b.t2 313.991
R3 b.t0 b.n11 41.3792
R4 b.n12 b.t0 40.2104
R5 b.n0 b.t6 28.5954
R6 b.n7 b.t8 28.5655
R7 b.n7 b.t5 28.5655
R8 b.n2 b.t1 28.5655
R9 b.n2 b.t12 28.5655
R10 b.n3 b.t14 28.5655
R11 b.n3 b.t10 28.5655
R12 b.n0 b.t4 26.3004
R13 b.n15 b.t7 26.2652
R14 b.n14 b.t9 26.2652
R15 b.n13 b.t13 26.2652
R16 b.n12 b.t11 26.2652
R17 b.n8 b.n7 25.3202
R18 b.n17 b.t15 13.2053
R19 b.n17 b.t3 6.63265
R20 b.n4 b.n2 1.62544
R21 b.n5 b.n4 1.44539
R22 b.n13 b.n12 0.718158
R23 b.n14 b.n13 0.718158
R24 b.n15 b.n14 0.718158
R25 b b.n18 0.594255
R26 b.n0 b.n15 0.517171
R27 b b.n16 0.502062
R28 b.n6 b.n5 0.191757
R29 b.n1 b.n6 0.189496
R30 b.n1 b.n10 0.162765
R31 b.n4 b.n3 0.156686
R32 b.n1 b.n0 0.0877146
R33 b.n10 b.n9 0.0870593
R34 b.n18 b.n17 0.0678366
R35 b.n16 b.n1 0.0614375
R36 b.n1 b.n8 0.0511368
R37 vd.n49 vd.n48 647.907
R38 vd.n49 vd.n32 647.529
R39 vd.t20 vd.t2 331.216
R40 vd.t2 vd.t17 331.216
R41 vd.t9 vd.t4 331.216
R42 vd.t6 vd.t9 331.216
R43 vd.t14 vd.t6 331.216
R44 vd.t41 vd.t35 331.216
R45 vd.t35 vd.t33 331.216
R46 vd.t33 vd.t29 331.216
R47 vd.t37 vd.t31 331.216
R48 vd.t23 vd.t37 331.216
R49 vd.n36 vd.t41 228.514
R50 vd.n35 vd.t14 210.542
R51 vd.t42 vd.t39 70.1694
R52 vd.t27 vd.t1 70.1694
R53 vd.t12 vd.t26 70.0291
R54 vd.t0 vd.t15 70.0291
R55 vd.n45 vd.t42 68.5376
R56 vd.t1 vd.n39 63.6434
R57 vd.n29 vd.t0 63.5148
R58 vd.t26 vd.n23 62.9732
R59 vd.n10 vd.t19 39.5312
R60 vd.n2 vd.t22 39.5292
R61 vd.n36 vd.n35 38.514
R62 vd.n42 vd.t27 37.5327
R63 vd.n26 vd.t12 35.2862
R64 vd.t15 vd.n26 34.7434
R65 vd.t39 vd.n42 32.6372
R66 vd.n2 vd.t25 28.6459
R67 vd.n0 vd.t36 28.5655
R68 vd.n0 vd.t34 28.5655
R69 vd.n1 vd.t38 28.5655
R70 vd.n1 vd.t24 28.5655
R71 vd.n4 vd.t30 28.5655
R72 vd.n4 vd.t32 28.5655
R73 vd.n11 vd.t21 28.5655
R74 vd.n11 vd.t3 28.5655
R75 vd.n13 vd.t18 28.5655
R76 vd.n13 vd.t5 28.5655
R77 vd.n30 vd.n29 21.216
R78 vd.n31 vd.n30 16.7426
R79 vd.n46 vd.t23 16.3842
R80 vd.n46 vd.n45 16.211
R81 vd.n30 vd.t20 12.5482
R82 vd.n47 vd.n46 7.64222
R83 vd.n21 vd.n9 5.78879
R84 vd.n8 vd.n7 5.72509
R85 vd.n19 vd.n18 2.24963
R86 vd.n7 vd.t40 1.90483
R87 vd.n7 vd.t28 1.90483
R88 vd.n9 vd.t13 1.90483
R89 vd.n9 vd.t16 1.90483
R90 vd.n8 vd.n6 1.79965
R91 vd.n14 vd.n12 1.56925
R92 vd.n5 vd.n3 1.5417
R93 vd.n15 vd.n14 1.438
R94 vd.n6 vd.n5 1.38515
R95 vd.n6 vd.n0 0.77517
R96 vd.n12 vd.n10 0.686006
R97 vd.n50 vd.n21 0.503104
R98 vd vd.n8 0.497524
R99 vd.n21 vd.n20 0.365502
R100 vd.n14 vd.n13 0.157684
R101 vd.n5 vd.n4 0.156686
R102 vd.n18 vd.n15 0.103522
R103 vd.n3 vd.n2 0.0791768
R104 vd.n18 vd.n17 0.0597867
R105 vd.n20 vd.n19 0.05675
R106 vd.n3 vd.n1 0.0493677
R107 vd.n12 vd.n11 0.0461626
R108 vd.n17 vd.n16 0.024973
R109 vd vd.n50 0.0239375
R110 vd.n25 vd.n24 0.00431884
R111 vd.n26 vd.n25 0.00431884
R112 vd.n41 vd.n40 0.00425193
R113 vd.n42 vd.n41 0.00425193
R114 vd.n48 vd.n47 0.00389051
R115 vd.n32 vd.n31 0.00389051
R116 vd.n44 vd.n43 0.0021559
R117 vd.n45 vd.n44 0.0021559
R118 vd.n28 vd.n27 0.00213065
R119 vd.n29 vd.n28 0.00213065
R120 vd.n39 vd.n38 0.00181202
R121 vd.n23 vd.n22 0.00181202
R122 vd.n34 vd.n33 0.0017783
R123 vd.n35 vd.n34 0.0017783
R124 vd.n49 vd.n37 0.000827345
R125 vd.n37 vd.n36 0.000827345
R126 vd.n50 vd.n49 0.000504092
R127 out.n4 out.t2 377.192
R128 out.n1 out.t0 377.175
R129 out.n7 out.t4 5.53268
R130 out.n6 out.t8 3.4805
R131 out.n6 out.t7 3.4805
R132 out.n7 out.n6 2.35238
R133 out.n5 out.n4 2.02858
R134 out.n2 out.n1 2.00736
R135 out.n3 out.t6 1.90483
R136 out.n3 out.t3 1.90483
R137 out.n0 out.t1 1.90483
R138 out.n0 out.t5 1.90483
R139 out.n8 out.n7 0.80675
R140 out out.n8 0.783312
R141 out.n8 out.n2 0.182565
R142 out.n7 out.n5 0.182565
R143 out.n5 out.n3 0.00195207
R144 out.n2 out.n0 0.00195207
R145 gnd.n23 gnd.n20 560.566
R146 gnd.n32 gnd.n27 547.013
R147 gnd.t21 gnd.t8 412.351
R148 gnd.t3 gnd.t10 412.351
R149 gnd.n30 gnd.t0 399.565
R150 gnd.n35 gnd.n32 374.579
R151 gnd.n21 gnd.t15 348.421
R152 gnd.t13 gnd.t3 263.712
R153 gnd.n41 gnd.n40 242.918
R154 gnd.n24 gnd.t21 217.363
R155 gnd.t0 gnd.n29 214.167
R156 gnd.n24 gnd.t5 194.988
R157 gnd.t2 gnd.t13 153.434
R158 gnd.n41 gnd.n23 147.294
R159 gnd.n33 gnd.t2 107.084
R160 gnd.t18 gnd.t4 107.084
R161 gnd.n13 gnd.t17 65.675
R162 gnd.n6 gnd.t14 65.5414
R163 gnd.n21 gnd.t23 63.9308
R164 gnd.n38 gnd.t18 35.1621
R165 gnd.n44 gnd.n43 31.16
R166 gnd.n43 gnd.t11 17.4005
R167 gnd.n43 gnd.t1 17.4005
R168 gnd.n40 gnd.n35 13.5534
R169 gnd.n30 gnd.t7 12.7866
R170 gnd.n38 gnd.t12 11.1883
R171 gnd.n13 gnd.t20 6.44128
R172 gnd.n44 gnd.n42 6.30056
R173 gnd.n42 gnd.n18 4.9255
R174 gnd.n7 gnd.t16 3.4805
R175 gnd.n7 gnd.t24 3.4805
R176 gnd.n14 gnd.t9 3.4805
R177 gnd.n14 gnd.t19 3.4805
R178 gnd.n0 gnd.t6 3.4805
R179 gnd.n0 gnd.t22 3.4805
R180 gnd.n8 gnd.n6 3.21916
R181 gnd.n15 gnd.n13 2.95318
R182 gnd gnd.n44 1.74425
R183 gnd.n9 gnd.n8 0.618
R184 gnd.n16 gnd.n15 0.60175
R185 gnd.n11 gnd.n5 0.412265
R186 gnd.n18 gnd.n16 0.139389
R187 gnd.n18 gnd.n17 0.139389
R188 gnd.n5 gnd.n3 0.0593235
R189 gnd.n32 gnd.n31 0.0431634
R190 gnd.n31 gnd.n30 0.0431634
R191 gnd.n23 gnd.n22 0.0388129
R192 gnd.n22 gnd.n21 0.0388129
R193 gnd.n11 gnd.n2 0.0285795
R194 gnd.n35 gnd.n34 0.0215341
R195 gnd.n34 gnd.n33 0.0215341
R196 gnd.n16 gnd.n12 0.01925
R197 gnd.n40 gnd.n39 0.00984699
R198 gnd.n39 gnd.n38 0.00984699
R199 gnd.n27 gnd.n26 0.007537
R200 gnd.n20 gnd.n19 0.007537
R201 gnd.n29 gnd.n28 0.00701261
R202 gnd.n41 gnd.n25 0.00701261
R203 gnd.n25 gnd.n24 0.00701261
R204 gnd.n37 gnd.n36 0.00517349
R205 gnd.n38 gnd.n37 0.00517349
R206 gnd.n12 gnd.n11 0.00425
R207 gnd.n11 gnd.n10 0.00425
R208 gnd.n10 gnd.n9 0.003
R209 gnd.n8 gnd.n7 0.00294771
R210 gnd.n15 gnd.n14 0.00294771
R211 gnd.n5 gnd.n4 0.00278445
R212 gnd.n1 gnd.n0 0.00193715
R213 gnd.n2 gnd.n1 0.00100999
R214 gnd.n42 gnd.n41 0.000506305
R215 d.n9 d.t1 377.216
R216 d.n8 d.t4 377.163
R217 d.n2 d.t13 134.298
R218 d.n4 d.t8 133.787
R219 d.n3 d.t6 133.761
R220 d.n2 d.t12 133.761
R221 d.n0 d.t3 5.55126
R222 d.n6 d.t7 3.4805
R223 d.n6 d.t9 3.4805
R224 d d.n7 3.10062
R225 d.n0 d.n9 2.02586
R226 d.n1 d.n8 1.99422
R227 d.n5 d.t0 1.91167
R228 d.n1 d.t11 1.90534
R229 d.n0 d.t10 1.90483
R230 d.n0 d.t2 1.90483
R231 d.n1 d.t5 1.89094
R232 d d.n1 0.77675
R233 d.n1 d.n0 0.647901
R234 d.n3 d.n2 0.538
R235 d.n4 d.n3 0.394346
R236 d.n7 d.n6 0.151643
R237 d.n5 d.n4 0.0558728
R238 d.n7 d.n5 0.0333947
R239 ib.n0 ib.t5 38.0465
R240 ib.n0 ib.t3 37.3602
R241 ib.n1 ib.t0 18.7496
R242 ib.n1 ib.t2 17.4934
R243 ib.n8 ib.t4 17.4005
R244 ib.n8 ib.t1 17.4005
R245 ib ib.n12 5.82847
R246 ib.n8 ib.n7 1.98351
R247 ib.n9 ib.n6 1.5912
R248 ib.n12 ib.n0 0.27692
R249 ib.n4 ib.n1 0.097375
R250 ib.n3 ib.n2 0.0963763
R251 ib.n11 ib.n10 0.0208125
R252 ib.n12 ib.n11 0.0174603
R253 ib.n4 ib.n3 0.0127549
R254 ib.n10 ib.n9 0.00846233
R255 ib.n9 ib.n8 0.00846233
R256 ib.n5 ib.n4 0.0051875
R257 ib.n10 ib.n5 0.003625
R258 in in.t0 325.817
C0 a vd 5.21f
C1 d vd 3.92f
C2 vd ib 0.0124f
C3 c out 0.0405f
C4 c b 0.16f
C5 in a 0.227f
C6 d in 0.673f
C7 in ib 0.573f
C8 a out 0.0961f
C9 d out 35.6f
C10 a b 0.239f
C11 d b 0.0351f
C12 out ib 0.0478f
C13 c a 0.199f
C14 in vd 0.376f
C15 d c 0.0518f
C16 c ib 0.185f
C17 vd out 4.72f
C18 b vd 6.07f
C19 d a 1.27f
C20 a ib 0.00973f
C21 c vd 0.00332f
C22 in out 0.0539f
C23 d ib 0.468f
C24 in b 0.112f
C25 b out 1.93f
C26 in c 0.416f
.ends

