** sch_path:
*+ /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/impedance-transformer_tb-ac2.sch
**.subckt impedance-transformer_tb-ac2
Vin1 net1 GND DC 0 AC 1
.save i(vin1)
R4 out net1 75 m=1
x2 out_ask out GND impedance-transformer
x1 vd out_ask GND GND ask-modulator
Vdd vd GND DC 1.8 AC 0
.save i(vdd)
**** begin user architecture code



.control
destroy all
save all
ac lin 1k 1k 4G
set units=degrees
run

set color0=white
set color1=black

plot smithgrid out
.endc

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


*C= 19.68521p R= 191.6

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/impedance-transformer.sym # of pins=3
** sym_path:
*+ /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/impedance-transformer.sym
** sch_path:
*+ /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/impedance-transformer.sch
.subckt impedance-transformer in out gnd
*.iopin gnd
*.iopin in
*.iopin out
XC0 in gnd sky130_fd_pr__cap_mim_m3_2 W=23.2 L=23.2 MF=9 m=9
XC1 out gnd sky130_fd_pr__cap_mim_m3_2 W=17.7 L=17.7 MF=25 m=25
x1 in out l1
**** begin user architecture code

* NGSPICE file created from impedance-transformer.ext - technology: sky





**** end user architecture code
.ends


* expanding   symbol:
*+  /home/hugodg/projects-sky130/temp-sensor/ask_modulator/xschem/ask-modulator.sym # of pins=4
** sym_path: /home/hugodg/projects-sky130/temp-sensor/ask_modulator/xschem/ask-modulator.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/ask_modulator/xschem/ask-modulator.sch
.subckt ask-modulator vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=24.4 L=24.4 MF=3 m=3
XR1 out vd gnd sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
x1 vd out l0
**** begin user architecture code


R0 vd vd.t1 0.714
R1 vd.t0 vd.t2 0.066
R2 vd.t1 vd.t0 0.066
R3 gnd.n15 gnd.n14 71.405
R4 gnd.n18 gnd.n17 71.152
R5 gnd.n6 gnd.n5 67.749
R6 gnd.n8 gnd.n7 67.387
R7 gnd gnd.n20 4.959
R8 gnd.n9 gnd.n8 1.449
R9 gnd.n20 gnd.n9 0.359
R10 gnd.n5 gnd.n4 0.13
R11 gnd.n20 gnd.n19 0.114
R12 gnd.n17 gnd.n16 0.109
R13 gnd.n19 gnd.n15 0.094
R14 gnd.n9 gnd.n6 0.031
R15 gnd.n11 gnd.n10 0.026
R16 gnd.n19 gnd.n18 0.017
R17 gnd.n12 gnd.n11 0.017
R18 gnd.n13 gnd.n12 0.01
R19 gnd.n2 gnd.n1 0.007
R20 gnd.n1 gnd.n0 0.007
R21 gnd.n3 gnd.n2 0.002
R22 gnd.n6 gnd.n3 0.001
R23 gnd.n15 gnd.n13 0.001
R24 in in.t0 396.948
C0 in gnd 0.07fF
C1 in out 0.25fF
C2 gnd vd 0.37fF
C3 vd out 3.12fF
C4 gnd out 0.33fF
C5 in 0 1.68fF
C6 vd.t2 0 36.61fF
C7 vd.t0 0 34.66fF
C8 vd.t1 0 49.33fF
C9 gnd 0 -0.63fF
C10 out 0 217.77fF
C11 vd 0 13.16fF


**** end user architecture code
XM1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/l1.sym
*+ # of pins=2
** sym_path: /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/l1.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/impedance-transformer/xschem/l1.sch
.subckt l1 p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 622.2p m=1
Cs1 p1 net1 57.26f m=1
Cs2 p2 net2 50.34f m=1
Rs1 net1 GND 17.57 m=1
Rs2 net2 GND 31.85 m=1
R1 p2 net3 2.202 m=1
.ends


* expanding   symbol:  /home/hugodg/projects-sky130/temp-sensor/ask_modulator/xschem/l0.sym # of
*+ pins=2
** sym_path: /home/hugodg/projects-sky130/temp-sensor/ask_modulator/xschem/l0.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/ask_modulator/xschem/l0.sch
.subckt l0 p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 993p m=1
Cs1 p1 net1 58.53f m=1
Cs2 p2 net2 52.93f m=1
Rs1 net1 GND 24.1 m=1
Rs2 net2 GND 22.94 m=1
R1 p2 net3 3.443 m=1
.ends

.GLOBAL GND
.end
