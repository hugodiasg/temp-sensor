magic
tech sky130A
magscale 1 2
timestamp 1700102200
<< nwell >>
rect -3160 2300 -2740 2540
rect -1049 2209 -840 2530
rect -400 2209 -260 2530
<< nsubdiff >>
rect -3060 2430 -2960 2450
rect -3060 2390 -3030 2430
rect -2990 2390 -2960 2430
rect -3060 2360 -2960 2390
<< nsubdiffcont >>
rect -3030 2390 -2990 2430
<< locali >>
rect -3060 2440 -2960 2450
rect -3060 2390 -3050 2440
rect -2980 2390 -2960 2440
rect -3060 2360 -2960 2390
<< viali >>
rect -3050 2430 -2980 2440
rect -3050 2390 -3030 2430
rect -3030 2390 -2990 2430
rect -2990 2390 -2980 2430
rect -120 2320 -80 2880
rect -2860 2160 -2820 2220
rect -830 2160 -790 2200
rect -2580 2090 -2520 2130
rect -1140 2040 -1080 2100
rect -120 1620 -80 1780
<< metal1 >>
rect -2940 4820 -2720 5220
rect -2580 4820 -2360 5220
rect -2260 4820 -2040 5220
rect -1920 4820 -1700 5220
rect -1440 4820 -1220 5220
rect -1100 4820 -880 5220
rect -780 4820 -560 5220
rect -440 4820 -220 5220
rect -140 5160 60 5360
rect -140 5000 -20 5160
rect -140 4920 -120 5000
rect -20 4920 -10 5000
rect -2980 3820 -2860 3900
rect -3180 3620 -2860 3820
rect -2980 3480 -2860 3620
rect -2760 3480 -2540 3880
rect -2420 3480 -2200 3880
rect -2100 3480 -1880 3880
rect -1740 3860 -1400 3880
rect -1740 3500 -1620 3860
rect -1540 3500 -1400 3860
rect -1740 3480 -1400 3500
rect -1260 3480 -1040 3880
rect -940 3480 -720 3880
rect -620 3480 -400 3880
rect -300 3440 -220 3520
rect -720 3420 -220 3440
rect -720 3360 -700 3420
rect -620 3360 -220 3420
rect -310 3280 -300 3300
rect -1630 3200 -1620 3280
rect -1540 3200 -300 3280
rect -220 3200 -210 3300
rect -1620 3180 -220 3200
rect -310 2940 -300 3000
rect -240 2980 -230 3000
rect -240 2940 -220 2980
rect -3180 2850 -2980 2920
rect -3180 2740 -580 2850
rect -510 2740 -500 2850
rect -3180 2720 -2980 2740
rect -3180 2540 -2980 2600
rect -3180 2440 -2840 2540
rect -3180 2400 -3050 2440
rect -3060 2390 -3050 2400
rect -2980 2390 -2960 2440
rect -3060 2360 -2960 2390
rect -410 2320 -400 2900
rect -340 2320 -300 2900
rect -126 2880 -74 2892
rect -220 2320 -120 2880
rect -80 2860 -40 2880
rect -40 2780 -30 2860
rect -80 2740 -40 2780
rect -40 2660 -30 2740
rect -80 2600 -40 2660
rect -40 2520 -30 2600
rect -80 2460 -40 2520
rect -40 2380 -30 2460
rect -80 2320 -40 2380
rect -126 2308 -74 2320
rect -3180 2220 -2980 2260
rect -2866 2220 -2814 2232
rect -3180 2160 -2860 2220
rect -2820 2160 -2814 2220
rect -3180 2060 -2980 2160
rect -2866 2148 -2814 2160
rect -842 2200 -778 2206
rect -590 2200 -580 2220
rect -842 2160 -830 2200
rect -790 2160 -580 2200
rect -842 2154 -778 2160
rect -590 2140 -580 2160
rect -500 2140 -490 2220
rect -300 2200 -280 2240
rect -290 2180 -280 2200
rect -220 2180 -210 2240
rect -2600 2070 -2590 2140
rect -2510 2070 -2500 2140
rect -2150 2080 -2140 2140
rect -2080 2080 -2070 2140
rect -1152 2100 -1068 2106
rect -1152 2040 -1140 2100
rect -1080 2040 -700 2100
rect -620 2040 -610 2100
rect -1152 2034 -1068 2040
rect -2870 1900 -2860 1980
rect -2780 1900 -2770 1980
rect -290 1900 -280 1920
rect -300 1860 -280 1900
rect -220 1860 -210 1920
rect -2590 1800 -2580 1860
rect -2520 1850 -350 1860
rect -2520 1800 -420 1850
rect -430 1790 -420 1800
rect -360 1800 -350 1850
rect -360 1790 -300 1800
rect -3180 1640 -2980 1700
rect -3180 1580 -2140 1640
rect -2080 1580 -2070 1640
rect -410 1620 -300 1790
rect -220 1780 -20 1800
rect -220 1760 -120 1780
rect -80 1760 -20 1780
rect -220 1620 -160 1760
rect -60 1620 -20 1760
rect -140 1600 -20 1620
rect -3180 1500 -2980 1580
rect -300 1540 -220 1580
rect -1760 -360 -1560 -320
rect -2900 -500 -2880 -360
rect -2780 -380 -60 -360
rect -2780 -500 -160 -380
rect -60 -500 -50 -380
rect -2900 -520 -60 -500
<< via1 >>
rect -120 4920 -20 5000
rect -1620 3500 -1540 3860
rect -700 3360 -620 3420
rect -1620 3200 -1540 3280
rect -300 3200 -220 3300
rect -300 2940 -240 3000
rect -580 2740 -510 2850
rect -400 2320 -340 2900
rect -120 2780 -80 2860
rect -80 2780 -40 2860
rect -120 2660 -80 2740
rect -80 2660 -40 2740
rect -120 2520 -80 2600
rect -80 2520 -40 2600
rect -120 2380 -80 2460
rect -80 2380 -40 2460
rect -580 2140 -500 2220
rect -280 2180 -220 2240
rect -2590 2130 -2510 2140
rect -2590 2090 -2580 2130
rect -2580 2090 -2520 2130
rect -2520 2090 -2510 2130
rect -2590 2070 -2510 2090
rect -2140 2080 -2080 2140
rect -700 2040 -620 2100
rect -2860 1900 -2780 1980
rect -280 1860 -220 1920
rect -2580 1800 -2520 1860
rect -420 1790 -360 1850
rect -2140 1580 -2080 1640
rect -160 1620 -120 1760
rect -120 1620 -80 1760
rect -80 1620 -60 1760
rect -2880 -500 -2780 -360
rect -160 -500 -60 -380
<< metal2 >>
rect -120 5000 -20 5010
rect -140 4920 -120 5000
rect -1620 3860 -1520 3880
rect -1540 3500 -1520 3860
rect -1620 3280 -1520 3500
rect -1540 3200 -1520 3280
rect -1620 3160 -1520 3200
rect -700 3420 -620 3430
rect -2590 2140 -2510 2150
rect -2590 2060 -2510 2070
rect -2140 2140 -2080 2150
rect -2860 1980 -2780 1990
rect -2880 1900 -2860 1980
rect -2880 -360 -2780 1900
rect -2580 1870 -2540 2060
rect -2580 1860 -2520 1870
rect -2580 1790 -2520 1800
rect -2140 1640 -2080 2080
rect -700 2100 -620 3360
rect -300 3300 -180 3310
rect -300 3170 -180 3180
rect -300 3000 -220 3170
rect -240 2940 -220 3000
rect -300 2930 -240 2940
rect -400 2900 -340 2910
rect -580 2850 -510 2860
rect -580 2230 -510 2740
rect -140 2860 -20 4920
rect -140 2780 -120 2860
rect -40 2780 -20 2860
rect -140 2740 -20 2780
rect -140 2660 -120 2740
rect -40 2660 -20 2740
rect -140 2600 -20 2660
rect -140 2520 -120 2600
rect -40 2520 -20 2600
rect -140 2460 -20 2520
rect -140 2380 -120 2460
rect -40 2380 -20 2460
rect -140 2320 -20 2380
rect -580 2220 -500 2230
rect -580 2130 -500 2140
rect -700 2030 -620 2040
rect -400 1860 -340 2320
rect -420 1850 -340 1860
rect -280 2240 -220 2250
rect -280 1920 -220 2180
rect -280 1850 -220 1860
rect -360 1790 -340 1850
rect -420 1780 -340 1790
rect -400 1620 -340 1780
rect -160 1760 -60 1780
rect -2140 1570 -2080 1580
rect -2880 -510 -2780 -500
rect -160 -380 -60 1620
rect -160 -510 -60 -500
<< via2 >>
rect -300 3200 -220 3300
rect -220 3200 -180 3300
rect -300 3180 -180 3200
rect -160 -480 -60 -380
<< metal3 >>
rect -320 3300 -160 3320
rect -320 3180 -300 3300
rect -180 3180 -160 3300
rect -320 3160 -160 3180
rect -180 -380 -40 -360
rect -200 -480 -160 -380
rect -60 -480 -40 -380
rect -200 -500 -40 -480
<< via3 >>
rect -300 3180 -180 3300
rect -160 -480 -60 -380
<< metal4 >>
rect -301 3300 -179 3301
rect -301 3180 -300 3300
rect -180 3180 440 3300
rect -301 3179 -179 3180
rect -180 -380 600 -360
rect -180 -480 -160 -380
rect -60 -480 600 -380
rect -161 -481 -59 -480
use sky130_fd_pr__res_xhigh_po_0p35_XMXTTL  sky130_fd_pr__res_xhigh_po_0p35_XMXTTL_0
timestamp 1700079212
transform 1 0 -840 0 1 4350
box -616 -882 616 882
use sky130_fd_pr__res_xhigh_po_0p35_XMXTTL  sky130_fd_pr__res_xhigh_po_0p35_XMXTTL_1
timestamp 1700079212
transform 1 0 -2314 0 1 4350
box -616 -882 616 882
use sky130_fd_sc_hd__dfrbp_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 -2882 0 1 1948
box -38 -48 2154 592
use sky130_fd_pr__cap_mim_m3_1_A4KLY5  XC1
timestamp 1700078798
transform 0 1 3000 -1 0 2426
box -2906 -2760 2906 2760
use sky130_fd_pr__nfet_01v8_648S5X  XN1
timestamp 1700078798
transform 1 0 -255 0 1 1714
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGSNAL  XP1
timestamp 1700078798
transform 1 0 -255 0 1 2593
box -211 -519 211 519
<< labels >>
flabel metal1 -3180 3620 -2980 3820 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal1 -3180 2060 -2980 2260 0 FreeSans 256 0 0 0 clk
port 2 nsew
flabel metal1 -3180 1500 -2980 1700 0 FreeSans 256 0 0 0 reset_b_dff
port 4 nsew
flabel metal1 -1760 -520 -1560 -320 0 FreeSans 256 0 0 0 gnd
port 1 nsew
flabel metal1 -3180 2720 -2980 2920 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 -140 5160 60 5360 0 FreeSans 256 0 0 0 vd
port 6 nsew
flabel metal1 -3180 2400 -2980 2600 0 FreeSans 256 0 0 0 vpwr
port 5 nsew
<< end >>
