magic
tech sky130B
timestamp 1644922882
<< metal1 >>
rect 3170 -870 4680 -820
rect 3170 -1050 3190 -870
rect 3550 -1050 4680 -870
rect 3170 -1090 4680 -1050
rect 5180 -860 6300 -810
rect 5180 -1040 5920 -860
rect 6280 -1040 6300 -860
rect 5180 -1080 6300 -1040
rect 4240 -1400 4340 -1090
rect 4430 -1290 5180 -1120
rect 4980 -1400 5180 -1290
rect 4240 -1420 4880 -1400
rect 3170 -1520 4880 -1420
rect 4240 -2250 4880 -1520
rect 4940 -1680 5180 -1400
rect 4940 -1870 5330 -1680
rect 4940 -2250 5180 -1870
rect 4860 -2580 4940 -2270
rect 3170 -2680 4940 -2580
rect 5240 -2990 5330 -1870
rect 3170 -3090 5330 -2990
rect 5480 -3340 5560 -1080
rect 3170 -3440 5560 -3340
<< via1 >>
rect 3190 -1050 3550 -870
rect 5920 -1040 6280 -860
<< metal2 >>
rect 3170 -870 3570 -850
rect 3170 -1050 3190 -870
rect 3550 -1050 3570 -870
rect 3170 -1090 3570 -1050
rect 5900 -860 6300 -840
rect 5900 -1040 5920 -860
rect 6280 -1040 6300 -860
rect 5900 -1080 6300 -1040
<< via2 >>
rect 3190 -1050 3550 -870
rect 5920 -1040 6280 -860
<< metal3 >>
rect 3170 -870 3570 -850
rect 3170 -1050 3190 -870
rect 3550 -1050 3570 -870
rect 3170 -1090 3570 -1050
rect 5900 -860 6300 -840
rect 5900 -1040 5920 -860
rect 6280 -1040 6300 -860
rect 5900 -1080 6300 -1040
<< via3 >>
rect 3190 -1050 3550 -870
rect 5920 -1040 6280 -860
<< metal4 >>
rect 3170 7400 6750 7800
rect 3170 -870 3570 7400
rect 4720 6860 5210 7400
rect 3170 -1050 3190 -870
rect 3550 -1050 3570 -870
rect 3170 -1090 3570 -1050
rect 5900 -860 6300 -840
rect 5900 -1040 5920 -860
rect 6280 -1040 6300 -860
rect 5900 -1080 6300 -1040
<< via4 >>
rect 8040 7330 8560 7870
rect 5920 -1040 6280 -860
<< metal5 >>
rect 8028 7870 8572 7882
rect 8028 7330 8040 7870
rect 8560 7330 8572 7870
rect 8028 7318 8572 7330
rect 4750 195 5150 200
rect 4750 -530 5168 195
rect 4750 -770 6300 -530
rect 5900 -860 6300 -770
rect 5900 -1040 5920 -860
rect 6280 -1040 6300 -860
rect 5900 -5580 6300 -1040
rect 5900 -6190 7120 -5580
use sky130_fd_pr__nfet_g5v0d10v5_ML7W5H  XM1
timestamp 1644922882
transform -1 0 4909 0 1 -1816
box -139 -564 139 564
use sky130_fd_pr__res_xhigh_po_0p35_NVRUDW  XR1
timestamp 1644922882
transform 0 1 4929 -1 0 -1050
box -101 -549 100 549
use l0  l0_0
timestamp 1644768986
transform 1 0 7100 0 -1 8800
box -600 0 15000 15000
use sky130_fd_pr__cap_mim_m3_2_EZRVX8  sky130_fd_pr__cap_mim_m3_2_EZRVX8_0
timestamp 1644922882
transform -1 0 4965 0 1 3530
box -1255 -3720 1265 3720
<< labels >>
flabel metal1 3170 -3440 3270 -3340 0 FreeSans 64 0 0 0 vd
port 3 nsew
flabel metal1 3170 -3090 3270 -2990 0 FreeSans 64 0 0 0 gnd
port 0 nsew
flabel metal1 3170 -2680 3270 -2580 0 FreeSans 64 0 0 0 in
port 1 nsew
flabel metal1 3170 -1520 3270 -1420 0 FreeSans 64 0 0 0 out
port 2 nsew
<< end >>
