** sch_path: /foss/designs/temp-sensor/device-complete/xschem/device-complete-tb.sch
**.subckt device-complete-tb
vpwr vpwr GND 1.8
V3 clk GND pulse 0 1.8 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 '
vdd vd GND 1.8
ibias vd ib 20u
VSS vs GND 0
x1 vd clk out vpwr ib GND out_buff out_sigma vts device-complete-pex
**** begin user architecture code

*cmd step stop

.save
.control
destroy all
save all
set color0=white
set color1=black
set temp=35
set hcopypscolor = 1
set wr_singlescale
option numdgt=7
tran 40p 10u
*let pot=-i(vdd)*vd
save all

plot vts out_sigma out_buff avg(out_buff)
plot out


*meas tran pot_avg avg pot from=0 to=5u
*plot pot pot_avg pot_rms

wrdata /foss/designs/temp-sensor/data/tran35.txt vts out_sigma out_buff out

*linearize out
*fft out
*hardcopy ~/fft56.ps mag(out_ask) xlimit 1G 4G ylimit 0 55u
*plot mag(out) xlimit 1G 4G ylimit 0 65u

*wrdata ./fft10.txt mag(out)




.endc



 .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/temp-sensor/device-complete/xschem/device-complete-pex.sym # of
*+ pins=9
** sym_path: /foss/designs/temp-sensor/device-complete/xschem/device-complete-pex.sym
** sch_path: /foss/designs/temp-sensor/device-complete/xschem/device-complete-pex.sch
.subckt device-complete-pex vd clk out vpwr ib gnd out_buff out_sigma vts
*.iopin vd
*.ipin clk
*.opin out
*.iopin vpwr
*.iopin ib
*.iopin gnd
*.opin vts
*.opin out_buff
*.opin out_sigma
**** begin user architecture code


* NGSPICE file created from device-complete.ext - technology: sky130A

*.subckt device-complete gnd clk out_sigma vts ib out_buff vd out vpwr
X0 gnd.t82 gnd.t79 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=1
X1 a_16688_5320# a_16854_3988# gnd.t36 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X2 buffer_0.a.t6 buffer_0.a.t4 buffer_0.a.t5 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0
+ ps=0 w=1.5 l=0.15
X3 sensor_0.a.t7 sensor_0.b.t20 gnd.t91 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X4 sensor_0.b.t15 sensor_0.b.t14 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X5 vd.t71 buffer_0.b.t16 out_buff.t8 vd.t70 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3
+ w=15 l=1
X6 a_15868_2881# a_14791_2515# a_15706_2515# vpwr.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69
+ as=0.0588 ps=0.7 w=0.42 l=0.15
X7 gnd.t97 vpwr.t30 a_15403_2515# gnd.t96 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63
+ w=0.42 l=0.15
X8 a_15546_5320# a_15712_3988# gnd.t42 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X9 vd.t16 buffer_0.a.t9 buffer_0.a.t10 vd.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X10 gnd.t115 sensor_0.b.t21 vtd.t7 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X11 a_15141_2515# a_14791_2515# a_15046_2515# vpwr.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765
+ as=0.0651 ps=0.73 w=0.42 l=0.15
X12 sensor_0.c sensor_0.c sensor_0.c vd.t41 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6
+ w=2 l=1
X13 buffer_0.d.t6 buffer_0.d.t4 buffer_0.d.t5 vd.t40 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0
+ ps=0 w=15 l=1
X14 gnd.t26 ib.t3 ib.t4 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X15 gnd.t78 gnd.t76 gnd.t77 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X16 a_14550_5320# a_14716_3988# gnd.t103 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X17 ib.t2 ib.t0 ib.t1 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X18 a_15815_2515# a_14625_2515# a_15706_2515# gnd.t107 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75
+ as=0.0711 ps=0.755 w=0.36 l=0.15
X19 vts.t16 vtd.t12 vtd.t13 vts.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 gnd.t35 sensor_0.b.t12 sensor_0.b.t13 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X21 a_16356_5320# a_16522_3988# gnd.t121 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X22 vtd.t9 vtd.t8 vts.t14 vts.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 gnd.t75 gnd.t73 gnd.t74 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X24 gnd.t29 sensor_0.b.t22 sensor_0.a.t6 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X25 gnd.t72 gnd.t70 gnd.t71 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X26 vtd.t6 sensor_0.b.t23 gnd.t30 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X27 out_sigma.t1 a_16445_2515# vpwr.t11 vpwr.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52
+ as=0.154 ps=1.34 w=1 l=0.15
X28 vts.t12 vtd.t22 vtd.t23 vts.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 buffer_0.b.t6 buffer_0.b.t5 vd.t69 vd.t68 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X30 vtd.t5 sensor_0.b.t24 gnd.t39 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X31 vpwr.t13 clk.t0 a_14625_2515# vpwr.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166
+ ps=1.8 w=0.64 l=0.15
X32 a_17020_5320# sigma-delta_0.x1.Q gnd.t128 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X33 vtd.t17 vtd.t16 vts.t10 vts.t9 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 vd.t67 buffer_0.b.t3 buffer_0.b.t4 vd.t66 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X35 a_15237_2515# a_14791_2515# a_15141_2515# gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1
+ as=0.0594 ps=0.69 w=0.36 l=0.15
X36 a_15706_2515# a_14625_2515# a_15359_2757# vpwr.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7
+ as=0.129 ps=1.18 w=0.42 l=0.15
X37 vd.t46 a_6126_29386# gnd.t98 sky130_fd_pr__res_xhigh_po_0p35 l=5
X38 sensor_0.b.t19 vtd.t24 sensor_0.c vd.t72 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58
+ w=2 l=1
X39 a_15359_2757# a_15141_2515# vpwr.t7 vpwr.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18
+ as=0.218 ps=2.2 w=0.84 l=0.15
X40 gnd.t88 clk.t1 a_14625_2515# gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36
+ w=0.42 l=0.15
X41 vts.t8 vtd.t14 vtd.t15 vts.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X42 vd.t65 buffer_0.b.t14 buffer_0.b.t15 vd.t64 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X43 gnd.t49 sensor_0.b.t10 sensor_0.b.t11 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X44 vpwr.t15 a_15706_2515# a_15881_2489# vpwr.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67
+ as=0.0567 ps=0.69 w=0.42 l=0.15
X45 buffer_0.a.t3 buffer_0.a.t2 buffer_0.a.t3 vd.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0
+ ps=0 w=1 l=1
X46 a_15046_2515# sigma-delta_0.x1.D vpwr.t21 vpwr.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73
+ as=0.109 ps=1.36 w=0.42 l=0.15
X47 vd.t56 sensor_0.a.t10 sensor_0.a.t11 vd.t55 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58
+ ps=4.58 w=2 l=1
X48 buffer_0.a.t12 buffer_0.a.t11 vd.t13 vd.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X49 a_15881_2489# a_15706_2515# a_16060_2515# gnd.t93 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36
+ as=0.064 ps=0.725 w=0.42 l=0.15
X50 buffer_0.b.t0 vts.t25 buffer_0.c gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248
+ ps=1.83 w=1.5 l=0.15
X51 sensor_0.b.t9 sensor_0.b.t8 gnd.t27 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X52 a_14882_5320# a_15048_3988# gnd.t90 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X53 gnd.t114 sensor_0.b.t25 sensor_0.a.t5 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X54 sigma-delta_0.x1.Q a_15881_2489# gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169
+ ps=1.82 w=0.65 l=0.15
X55 vts.t24 vts.t21 vts.t23 vts.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X56 buffer_0.d.t1 buffer_0.a.t16 vd.t11 vd.t10 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17
+ ps=15.3 w=15 l=1
X57 out_buff.t10 buffer_0.d.t11 sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X58 a_15359_2757# a_15141_2515# gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135
+ ps=1.15 w=0.64 l=0.15
X59 vpwr.t29 a_15359_2757# a_15249_2881# vpwr.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755
+ as=0.116 ps=0.97 w=0.42 l=0.15
X60 a_15706_2515# a_14791_2515# a_15359_2757# gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755
+ as=0.0999 ps=0.985 w=0.36 l=0.15
X61 gnd.t83 sensor_0.b.t26 vtd.t4 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X62 vd.t37 vtd.t25 vts.t4 vd.t36 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X63 a_15214_5320# a_15380_3988# gnd.t48 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X64 vd.t35 vd.t32 vd.t34 vd.t33 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X65 gnd.t69 gnd.t67 gnd.t68 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X66 sensor_0.c vtd.t26 sensor_0.b.t17 vd.t39 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29
+ w=2 l=1
X67 out_buff.t5 out_buff.t3 out_buff.t4 vd.t43 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0
+ w=15 l=1
X68 out_sigma.t0 a_16445_2515# gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1
+ ps=0.985 w=0.65 l=0.15
X69 vd.t31 vd.t28 vd.t30 vd.t29 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X70 sensor_0.a.t4 sensor_0.b.t27 gnd.t31 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X71 sensor_0.a.t3 sensor_0.b.t28 gnd.t110 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X72 sigma-delta_0.x1.Q a_15881_2489# vpwr.t5 vpwr.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56
+ as=0.213 ps=1.67 w=1 l=0.15
X73 sensor_0.a.t9 sensor_0.a.t8 vd.t54 vd.t53 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29
+ ps=2.29 w=2 l=1
X74 vd.t73 out.t3 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X75 a_16060_2515# vpwr.t31 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125
+ ps=1.01 w=0.42 l=0.15
X76 gnd.t38 buffer_0.d.t12 out_buff.t0 gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725
+ ps=5.29 w=5 l=1
X77 buffer_0.c out_buff.t11 buffer_0.a.t15 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83
+ as=0.248 ps=1.83 w=1.5 l=0.15
X78 a_16024_5320# a_16190_3988# gnd.t108 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X79 out_buff.t7 buffer_0.d.t13 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725
+ ps=5.29 w=5 l=1
X80 sensor_0.b.t7 sensor_0.b.t6 gnd.t28 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X81 vd.t27 vd.t25 vd.t27 vd.t26 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X82 gnd.t22 sensor_0.b.t29 vtd.t3 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X83 gnd.t86 buffer_0.d.t9 buffer_0.d.t10 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725
+ ps=5.29 w=5 l=1
X84 a_16688_5320# a_16522_3988# gnd.t47 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X85 vd.t24 vd.t21 vd.t23 vd.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X86 vd.t63 buffer_0.b.t7 buffer_0.b.t8 vd.t62 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X87 buffer_0.d.t8 buffer_0.d.t7 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725
+ ps=5.29 w=5 l=1
X88 sensor_0.c sensor_0.a.t12 sensor_0.d vd.t52 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29
+ ps=2.29 w=2 l=1
X89 sensor_0.d sensor_0.a.t13 sensor_0.c vd.t51 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58
+ ps=4.58 w=2 l=1
X90 a_15546_5320# a_15380_3988# gnd.t89 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X91 buffer_0.d.t3 buffer_0.d.t2 buffer_0.d.t3 vd.t47 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0
+ ps=0 w=15 l=1
X92 vpwr.t3 a_15881_2489# a_15868_2881# vpwr.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81
+ as=0.0567 ps=0.69 w=0.42 l=0.15
X93 gnd.t66 gnd.t64 gnd.t65 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X94 gnd.t63 gnd.t61 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=1
X95 gnd.t60 gnd.t58 gnd.t59 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X96 gnd.t57 gnd.t54 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X97 buffer_0.c buffer_0.c buffer_0.c gnd.t113 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=1.08
+ ps=8.82 w=1 l=1
X98 vd.t20 vd.t17 vd.t19 vd.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X99 a_15046_2515# sigma-delta_0.x1.D gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745
+ as=0.221 ps=1.89 w=0.42 l=0.15
X100 vtd.t11 vtd.t10 vts.t6 vts.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X101 vd.t9 buffer_0.a.t17 buffer_0.d.t0 vd.t8 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17
+ ps=15.3 w=15 l=1
X102 gnd.t10 sensor_0.b.t4 sensor_0.b.t5 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X103 buffer_0.c ib.t5 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1
+ l=1
X104 vts.t3 vtd.t20 vtd.t21 vts.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X105 buffer_0.b.t13 buffer_0.b.t11 buffer_0.b.t12 vd.t61 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58
+ as=0 ps=0 w=1 l=1
X106 gnd.t8 sensor_0.b.t30 sensor_0.a.t2 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X107 a_15141_2515# a_14625_2515# a_15046_2515# gnd.t106 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69
+ as=0.066 ps=0.745 w=0.36 l=0.15
X108 vtd.t2 sensor_0.b.t31 gnd.t94 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X109 a_16356_5320# a_16190_3988# gnd.t92 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X110 vtd.t19 vtd.t18 vts.t1 vts.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X111 vtd.t1 sensor_0.b.t32 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X112 vd.t1 a_15712_3988# sigma-delta_0.x1.D vd.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87
+ ps=6.58 w=3 l=0.15
X113 sensor_0.c vtd.t27 sensor_0.b.t16 vd.t38 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29
+ ps=2.29 w=2 l=1
X114 a_15214_5320# a_15048_3988# gnd.t6 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X115 out_buff.t9 buffer_0.b.t17 vd.t60 vd.t59 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17
+ ps=15.3 w=15 l=1
X116 buffer_0.a.t8 buffer_0.a.t7 vd.t7 vd.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X117 vd.t74 out.t2 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X118 vd.t5 buffer_0.a.t13 buffer_0.a.t14 vd.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X119 sensor_0.b.t18 vtd.t28 sensor_0.c vd.t48 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29
+ ps=2.29 w=2 l=1
X120 a_17020_5320# a_16854_3988# gnd.t102 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X121 gnd.t116 sensor_0.b.t2 sensor_0.b.t3 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X122 sensor_0.d vtd.t29 vd.t45 vd.t44 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2
+ l=1
X123 a_14791_2515# a_14625_2515# vpwr.t18 vpwr.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8
+ as=0.0864 ps=0.91 w=0.64 l=0.15
X124 buffer_0.a.t1 buffer_0.a.t0 vd.t3 vd.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X125 a_14882_5320# a_14716_3988# gnd.t84 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X126 gnd.t14 a_15712_3988# sigma-delta_0.x1.D gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58
+ as=0.29 ps=2.58 w=1 l=0.15
X127 sensor_0.d sensor_0.a.t14 sensor_0.c vd.t50 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29
+ ps=2.29 w=2 l=1
X128 vts.t20 vts.t17 vts.t19 vts.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X129 a_14791_2515# a_14625_2515# gnd.t105 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36
+ as=0.0567 ps=0.69 w=0.42 l=0.15
X130 a_15249_2881# a_14625_2515# a_15141_2515# vpwr.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97
+ as=0.0724 ps=0.765 w=0.42 l=0.15
X131 buffer_0.b.t10 buffer_0.b.t9 buffer_0.b.t10 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83
+ as=0 ps=0 w=1.5 l=0.15
X132 sensor_0.b.t1 sensor_0.b.t0 gnd.t117 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X133 gnd.t109 sensor_0.b.t33 sensor_0.a.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X134 a_16024_5320# a_15712_3988# gnd.t125 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X135 vd.t75 out.t1 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X136 gnd.t112 out_sigma.t2 out.t0 gnd.t111 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ w=2 l=0.15
X137 sensor_0.c sensor_0.a.t15 sensor_0.d vd.t49 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29
+ ps=2.29 w=2 l=1
X138 gnd.t34 sensor_0.b.t34 vtd.t0 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X139 gnd.t3 a_15881_2489# a_15815_2515# gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669
+ ps=0.75 w=0.42 l=0.15
X140 a_15403_2515# a_15359_2757# a_15237_2515# gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63
+ as=0.14 ps=1.1 w=0.42 l=0.15
X141 a_15249_2881# vpwr.t25 vpwr.t27 vpwr.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703
+ ps=0.755 w=0.42 l=0.15
X142 a_15881_2489# vpwr.t22 vpwr.t24 vpwr.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69
+ as=0.0819 ps=0.81 w=0.42 l=0.15
X143 gnd.t1 a_15881_2489# a_16445_2515# gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109
+ ps=1.36 w=0.42 l=0.15
X144 a_14550_5320# out_buff.t6 gnd.t95 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X145 sensor_0.a.t0 sensor_0.b.t35 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X146 vpwr.t1 a_15881_2489# a_16445_2515# vpwr.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34
+ as=0.166 ps=1.8 w=0.64 l=0.15
X147 gnd.t53 gnd.t50 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X148 buffer_0.b.t2 buffer_0.b.t1 vd.t58 vd.t57 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X149 a_15712_3988# gnd.t12 sky130_fd_pr__cap_mim_m3_1 l=27.2 w=27.2
X150 out_buff.t2 out_buff.t1 out_buff.t2 vd.t42 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0
+ w=15 l=1
R0 gnd.n150 gnd.n3 16393.5
R1 gnd.n67 gnd.n61 9068.36
R2 gnd.n150 gnd.n149 4031.02
R3 gnd.n61 gnd.n60 1756.55
R4 gnd.n153 gnd.n150 1057.91
R5 gnd.n61 gnd.t128 905.341
R6 gnd.t125 gnd.t42 718.744
R7 gnd.n191 gnd.n190 585
R8 gnd.n245 gnd.n244 585
R9 gnd.n247 gnd.n246 585
R10 gnd.n2 gnd.n1 585
R11 gnd.n8 gnd.n5 560.566
R12 gnd.n142 gnd.n139 547.013
R13 gnd.n55 gnd.n54 523.47
R14 gnd.n26 gnd.t43 389.486
R15 gnd.t128 gnd.t102 382.409
R16 gnd.t102 gnd.t36 382.409
R17 gnd.t36 gnd.t47 382.409
R18 gnd.t47 gnd.t121 382.409
R19 gnd.t121 gnd.t92 382.409
R20 gnd.t92 gnd.t108 382.409
R21 gnd.t108 gnd.t125 382.409
R22 gnd.t42 gnd.t89 382.409
R23 gnd.t89 gnd.t48 382.409
R24 gnd.t48 gnd.t6 382.409
R25 gnd.t6 gnd.t90 382.409
R26 gnd.t90 gnd.t84 382.409
R27 gnd.t84 gnd.t103 382.409
R28 gnd.t103 gnd.t95 382.409
R29 gnd.n6 gnd.t62 348.421
R30 gnd.n155 gnd.t23 334.93
R31 gnd.n253 gnd.t7 331.329
R32 gnd.t11 gnd.t122 305.267
R33 gnd.t9 gnd.n192 298.916
R34 gnd.t124 gnd.t113 263.712
R35 gnd.n193 gnd.t19 262.902
R36 gnd.n146 gnd.n145 256.471
R37 gnd.n54 gnd.n53 247.828
R38 gnd.n134 gnd.n129 242.918
R39 gnd.n221 gnd.t21 223.286
R40 gnd.n127 gnd.t85 217.363
R41 gnd.n80 gnd.t120 215.036
R42 gnd.n143 gnd.t25 214.167
R43 gnd.t119 gnd.t104 211.339
R44 gnd.n143 gnd.t40 198.185
R45 gnd.n127 gnd.t99 194.988
R46 gnd.t95 gnd.n33 193.508
R47 gnd.t55 gnd.n154 172.868
R48 gnd.n223 gnd.n220 163.766
R49 gnd.t0 gnd.t4 159.876
R50 gnd.t4 gnd.t93 159.876
R51 gnd.n255 gnd.n245 156.236
R52 gnd.n90 gnd.t5 154.317
R53 gnd.n202 gnd.n201 153.976
R54 gnd.t118 gnd.t124 153.434
R55 gnd.n154 gnd.n153 152.16
R56 gnd.n200 gnd.n195 150.648
R57 gnd.n202 gnd.n191 148.707
R58 gnd.n129 gnd.n8 147.294
R59 gnd.t126 gnd.t33 141.167
R60 gnd.t13 gnd.n26 134.364
R61 gnd.n145 gnd.n142 133.742
R62 gnd.n92 gnd.n91 128.757
R63 gnd.t51 gnd.n252 127.85
R64 gnd.t45 gnd.t2 126.71
R65 gnd.n221 gnd.t17 118.847
R66 gnd.n88 gnd.n87 116.754
R67 gnd.t15 gnd.t96 112.254
R68 gnd.n252 gnd.n251 110.743
R69 gnd.n119 gnd.n78 107.24
R70 gnd.n106 gnd.n84 107.24
R71 gnd.t80 gnd.t11 107.084
R72 gnd.n23 gnd.n22 104.427
R73 gnd.n87 gnd.t46 100.001
R74 gnd.n31 gnd.n30 98.6358
R75 gnd.t107 gnd.t32 92.6947
R76 gnd.n149 gnd.n148 86.3064
R77 gnd.t32 gnd.t15 84.1907
R78 gnd.t43 gnd.t0 82.4899
R79 gnd.t2 gnd.t107 81.6395
R80 gnd.t33 gnd.t106 81.6395
R81 gnd.t106 gnd.t119 80.7891
R82 gnd.n193 gnd.t9 79.2311
R83 gnd.t93 gnd.t45 77.3874
R84 gnd.n84 gnd.t97 72.8576
R85 gnd.n87 gnd.t3 70.0005
R86 gnd.t104 gnd.t87 69.6181
R87 gnd.n157 gnd.n2 65.8829
R88 gnd.n15 gnd.t79 65.675
R89 gnd.n9 gnd.t61 65.5414
R90 gnd.t7 gnd.n248 64.8256
R91 gnd.n6 gnd.t37 63.9308
R92 gnd.t96 gnd.t126 61.2297
R93 gnd.n84 gnd.t16 60.5809
R94 gnd.n91 gnd.t1 57.1434
R95 gnd.t87 gnd.n23 53.8718
R96 gnd.n255 gnd.n247 48.5652
R97 gnd.n78 gnd.t105 38.5719
R98 gnd.n78 gnd.t88 38.5719
R99 gnd.n237 gnd.t50 37.3602
R100 gnd.n240 gnd.t76 37.3602
R101 gnd.n243 gnd.t58 37.3602
R102 gnd.n162 gnd.t70 37.3602
R103 gnd.n165 gnd.t64 37.3602
R104 gnd.n168 gnd.t73 37.3602
R105 gnd.n132 gnd.t80 35.1621
R106 gnd.n108 gnd.n107 34.6358
R107 gnd.n108 gnd.n82 34.6358
R108 gnd.n112 gnd.n82 34.6358
R109 gnd.n113 gnd.n112 34.6358
R110 gnd.n114 gnd.n113 34.6358
R111 gnd.n100 gnd.n99 34.6358
R112 gnd.n101 gnd.n100 34.6358
R113 gnd.n101 gnd.n85 34.6358
R114 gnd.n105 gnd.n85 34.6358
R115 gnd.n95 gnd.n94 34.6358
R116 gnd.n96 gnd.n95 34.6358
R117 gnd.n118 gnd.n80 29.7417
R118 gnd.n94 gnd.n90 27.8593
R119 gnd.n91 gnd.t44 25.4291
R120 gnd.n53 gnd.t111 24.5503
R121 gnd.n120 gnd.n119 24.4919
R122 gnd.n44 gnd.n41 24.3682
R123 gnd.n199 gnd.n196 23.4095
R124 gnd.n60 gnd.t98 22.9965
R125 gnd.t98 gnd.n55 22.9965
R126 gnd.n119 gnd.n118 22.9652
R127 gnd.n149 gnd.t118 20.7778
R128 gnd.n159 gnd.t54 18.6812
R129 gnd.n234 gnd.t67 18.6809
R130 gnd.n96 gnd.n88 17.6946
R131 gnd.n217 gnd.t83 17.4089
R132 gnd.n187 gnd.t116 17.4089
R133 gnd.n228 gnd.t29 17.4084
R134 gnd.n226 gnd.t109 17.4084
R135 gnd.n225 gnd.t114 17.4084
R136 gnd.n228 gnd.t31 17.4084
R137 gnd.n226 gnd.t110 17.4084
R138 gnd.n225 gnd.t18 17.4084
R139 gnd.n217 gnd.t20 17.4079
R140 gnd.n187 gnd.t117 17.4079
R141 gnd.n230 gnd.t91 17.4074
R142 gnd.n230 gnd.t8 17.4074
R143 gnd.n204 gnd.t22 17.4069
R144 gnd.n204 gnd.t30 17.4055
R145 gnd.n233 gnd.t69 17.405
R146 gnd.n233 gnd.t68 17.405
R147 gnd.n236 gnd.t53 17.405
R148 gnd.n236 gnd.t52 17.405
R149 gnd.n239 gnd.t78 17.405
R150 gnd.n239 gnd.t77 17.405
R151 gnd.n242 gnd.t60 17.405
R152 gnd.n242 gnd.t59 17.405
R153 gnd.n158 gnd.t57 17.405
R154 gnd.n158 gnd.t56 17.405
R155 gnd.n161 gnd.t72 17.405
R156 gnd.n161 gnd.t71 17.405
R157 gnd.n164 gnd.t66 17.405
R158 gnd.n164 gnd.t65 17.405
R159 gnd.n167 gnd.t75 17.405
R160 gnd.n167 gnd.t74 17.405
R161 gnd.n21 gnd.t14 17.405
R162 gnd.n206 gnd.t94 17.4034
R163 gnd.n205 gnd.t115 17.4034
R164 gnd.n212 gnd.t39 17.4034
R165 gnd.n211 gnd.t34 17.4034
R166 gnd.n182 gnd.t27 17.4034
R167 gnd.n181 gnd.t49 17.4034
R168 gnd.n176 gnd.t28 17.4034
R169 gnd.n175 gnd.t10 17.4034
R170 gnd.n171 gnd.t24 17.4034
R171 gnd.n170 gnd.t35 17.4034
R172 gnd.n135 gnd.t41 17.4005
R173 gnd.n135 gnd.t26 17.4005
R174 gnd.n114 gnd.n80 14.6829
R175 gnd.n146 gnd.n134 13.5534
R176 gnd.n140 gnd.t127 12.7866
R177 gnd.n132 gnd.t101 11.1883
R178 gnd.n92 gnd.n90 10.9075
R179 gnd.n253 gnd.t51 10.8047
R180 gnd.n21 gnd.n20 9.33321
R181 gnd.n157 gnd.n156 9.3005
R182 gnd.n156 gnd.n155 9.3005
R183 gnd.n202 gnd.n194 9.3005
R184 gnd.n194 gnd.n193 9.3005
R185 gnd.n223 gnd.n222 9.3005
R186 gnd.n222 gnd.n221 9.3005
R187 gnd.n255 gnd.n254 9.3005
R188 gnd.n254 gnd.n253 9.3005
R189 gnd.n49 gnd.t112 8.70236
R190 gnd.n107 gnd.n106 7.90638
R191 gnd.n155 gnd.t55 7.20328
R192 gnd.n15 gnd.t82 6.44128
R193 gnd.n126 gnd.n125 5.41306
R194 gnd.n137 gnd.n136 5.41306
R195 gnd.n116 gnd.n80 4.6505
R196 gnd.n94 gnd.n93 4.6505
R197 gnd.n95 gnd.n89 4.6505
R198 gnd.n97 gnd.n96 4.6505
R199 gnd.n99 gnd.n98 4.6505
R200 gnd.n100 gnd.n86 4.6505
R201 gnd.n102 gnd.n101 4.6505
R202 gnd.n103 gnd.n85 4.6505
R203 gnd.n105 gnd.n104 4.6505
R204 gnd.n107 gnd.n83 4.6505
R205 gnd.n109 gnd.n108 4.6505
R206 gnd.n110 gnd.n82 4.6505
R207 gnd.n112 gnd.n111 4.6505
R208 gnd.n113 gnd.n81 4.6505
R209 gnd.n115 gnd.n114 4.6505
R210 gnd.n118 gnd.n117 4.6505
R211 gnd.n119 gnd.n79 4.6505
R212 gnd.n76 gnd.n75 4.5005
R213 gnd.n77 gnd.n75 4.5005
R214 gnd gnd.n123 3.79922
R215 gnd.n12 gnd.t100 3.4805
R216 gnd.n12 gnd.t86 3.4805
R217 gnd.n10 gnd.t63 3.4805
R218 gnd.n10 gnd.t38 3.4805
R219 gnd.n16 gnd.t123 3.4805
R220 gnd.n16 gnd.t81 3.4805
R221 gnd.n11 gnd.n9 3.21916
R222 gnd.n17 gnd.n15 2.95318
R223 gnd.n74 gnd.n73 2.6505
R224 gnd.n99 gnd.n88 2.63579
R225 gnd.n49 gnd 2.5773
R226 gnd.n125 gnd.n124 2.43634
R227 gnd.n121 gnd.n75 2.25328
R228 gnd gnd.n0 2.00418
R229 gnd.n106 gnd.n105 1.88285
R230 gnd.n74 gnd.t12 1.47915
R231 gnd.n137 gnd.n135 1.41862
R232 gnd.n124 gnd.n74 1.22706
R233 gnd gnd.n0 1.2022
R234 gnd.n23 gnd 0.928252
R235 gnd.n136 gnd 0.793114
R236 gnd.n259 gnd.n258 0.685777
R237 gnd.n14 gnd.n11 0.6455
R238 gnd.n18 gnd.n17 0.62925
R239 gnd.n68 gnd.n32 0.54125
R240 gnd.n32 gnd.n31 0.541165
R241 gnd.n210 gnd.n204 0.447415
R242 gnd.n216 gnd.n210 0.438
R243 gnd.n218 gnd.n216 0.438
R244 gnd.n126 gnd.n19 0.425505
R245 gnd.n180 gnd.n174 0.375501
R246 gnd.n219 gnd.n218 0.375501
R247 gnd.n186 gnd.n180 0.3755
R248 gnd.n188 gnd.n186 0.3755
R249 gnd.n227 gnd.n225 0.373217
R250 gnd.n229 gnd.n227 0.371401
R251 gnd.n231 gnd.n229 0.369555
R252 gnd.n52 gnd.n48 0.366293
R253 gnd.n39 gnd.n38 0.365897
R254 gnd.n53 gnd.n39 0.365897
R255 gnd.n48 gnd.n47 0.365897
R256 gnd.n66 gnd.n65 0.347558
R257 gnd.n65 gnd.n64 0.347269
R258 gnd.n232 gnd.n231 0.338503
R259 gnd.n189 gnd.n188 0.330858
R260 gnd.n189 gnd.n169 0.290469
R261 gnd.n219 gnd.n203 0.281539
R262 gnd.n224 gnd.n219 0.245825
R263 gnd.n257 gnd.n232 0.244548
R264 gnd.n259 gnd.n0 0.230614
R265 gnd.n232 gnd.n224 0.180349
R266 gnd.n203 gnd.n189 0.156539
R267 gnd.n93 gnd.n92 0.144332
R268 gnd.n35 gnd.n34 0.1305
R269 gnd.t98 gnd.n35 0.1305
R270 gnd.n57 gnd.n56 0.1305
R271 gnd.t98 gnd.n57 0.1305
R272 gnd.n93 gnd.n89 0.120292
R273 gnd.n97 gnd.n89 0.120292
R274 gnd.n98 gnd.n97 0.120292
R275 gnd.n98 gnd.n86 0.120292
R276 gnd.n102 gnd.n86 0.120292
R277 gnd.n103 gnd.n102 0.120292
R278 gnd.n104 gnd.n103 0.120292
R279 gnd.n104 gnd.n83 0.120292
R280 gnd.n109 gnd.n83 0.120292
R281 gnd.n110 gnd.n109 0.120292
R282 gnd.n111 gnd.n110 0.120292
R283 gnd.n111 gnd.n81 0.120292
R284 gnd.n115 gnd.n81 0.120292
R285 gnd.n116 gnd.n115 0.120292
R286 gnd.n117 gnd.n116 0.120292
R287 gnd.n117 gnd.n79 0.120292
R288 gnd.n28 gnd.n27 0.10956
R289 gnd.t13 gnd.n28 0.10956
R290 gnd.n29 gnd.t13 0.10956
R291 gnd.n30 gnd.n29 0.10956
R292 gnd.n43 gnd.n42 0.10956
R293 gnd.n46 gnd.n45 0.10956
R294 gnd.t111 gnd.n46 0.10956
R295 gnd.n44 gnd.n43 0.109135
R296 gnd.n66 gnd.n63 0.0849523
R297 gnd.n63 gnd.n62 0.0845034
R298 gnd.n260 gnd.n259 0.0772045
R299 gnd.n260 gnd 0.0755
R300 gnd.n79 gnd.n76 0.0734167
R301 gnd.n235 gnd.n234 0.073412
R302 gnd.n160 gnd.n159 0.0734113
R303 gnd.n19 gnd.n18 0.063
R304 gnd.n161 gnd.n160 0.0610469
R305 gnd.n162 gnd.n161 0.0610469
R306 gnd.n164 gnd.n163 0.0610469
R307 gnd.n165 gnd.n164 0.0610469
R308 gnd.n167 gnd.n166 0.0610469
R309 gnd.n168 gnd.n167 0.0610469
R310 gnd.n236 gnd.n235 0.0610469
R311 gnd.n237 gnd.n236 0.0610469
R312 gnd.n239 gnd.n238 0.0610469
R313 gnd.n240 gnd.n239 0.0610469
R314 gnd.n242 gnd.n241 0.0610469
R315 gnd.n243 gnd.n242 0.0610469
R316 gnd.n256 gnd.n243 0.0573558
R317 gnd.n169 gnd.n168 0.0573547
R318 gnd.n257 gnd.n256 0.0464211
R319 gnd.n142 gnd.n141 0.0431634
R320 gnd.n141 gnd.n140 0.0431634
R321 gnd.n163 gnd.n162 0.0426875
R322 gnd.n166 gnd.n165 0.0426875
R323 gnd.n238 gnd.n237 0.0426875
R324 gnd.n241 gnd.n240 0.0426875
R325 gnd.n25 gnd.n24 0.0425017
R326 gnd.n26 gnd.n25 0.0425017
R327 gnd.n258 gnd 0.0395625
R328 gnd.n8 gnd.n7 0.0388129
R329 gnd.n7 gnd.n6 0.0388129
R330 gnd gnd.n260 0.0345909
R331 gnd.n77 gnd 0.0330521
R332 gnd.n124 gnd 0.03175
R333 gnd.n159 gnd.n158 0.031274
R334 gnd.n234 gnd.n233 0.0312734
R335 gnd.n122 gnd.n76 0.0265417
R336 gnd.n41 gnd.n40 0.0264102
R337 gnd.n120 gnd 0.0226354
R338 gnd.n147 gnd.n146 0.0215341
R339 gnd.n148 gnd.n147 0.0215341
R340 gnd.n18 gnd.n14 0.01675
R341 gnd.n218 gnd.n217 0.0153409
R342 gnd.n215 gnd.n213 0.0129048
R343 gnd.n122 gnd.n121 0.0114272
R344 gnd.n209 gnd.n207 0.0114167
R345 gnd.n121 gnd.n120 0.0113582
R346 gnd.n123 gnd.n75 0.0110001
R347 gnd.n134 gnd.n133 0.00984699
R348 gnd.n133 gnd.n132 0.00984699
R349 gnd.n201 gnd.n200 0.0092427
R350 gnd.n200 gnd.n199 0.0092427
R351 gnd.n250 gnd.n249 0.00883856
R352 gnd.n251 gnd.n250 0.00883856
R353 gnd.n152 gnd.n151 0.00883856
R354 gnd.n153 gnd.n152 0.00883856
R355 gnd.n71 gnd.n21 0.00867757
R356 gnd.n188 gnd.n187 0.00792873
R357 gnd.n37 gnd.n36 0.00762598
R358 gnd.n55 gnd.n37 0.00762598
R359 gnd.n59 gnd.n58 0.00762598
R360 gnd.n60 gnd.n59 0.00762598
R361 gnd.n5 gnd.n4 0.007537
R362 gnd.n139 gnd.n138 0.007537
R363 gnd.n145 gnd.n144 0.00701261
R364 gnd.n144 gnd.n143 0.00701261
R365 gnd.n129 gnd.n128 0.00701261
R366 gnd.n128 gnd.n127 0.00701261
R367 gnd.n73 gnd.n71 0.00634112
R368 gnd gnd.n77 0.00570833
R369 gnd.n185 gnd.n183 0.00546432
R370 gnd.n131 gnd.n130 0.00517349
R371 gnd.n132 gnd.n131 0.00517349
R372 gnd.n172 gnd.n170 0.00502806
R373 gnd.n177 gnd.n175 0.00502806
R374 gnd.n183 gnd.n181 0.00502805
R375 gnd.n207 gnd.n205 0.00502803
R376 gnd.n213 gnd.n211 0.00502803
R377 gnd.n198 gnd.n197 0.00487141
R378 gnd.n199 gnd.n198 0.00487141
R379 gnd.n69 gnd.n68 0.00441022
R380 gnd.n172 gnd.n171 0.00402807
R381 gnd.n177 gnd.n176 0.00402806
R382 gnd.n183 gnd.n182 0.00402806
R383 gnd.n207 gnd.n206 0.00402804
R384 gnd.n213 gnd.n212 0.00402803
R385 gnd.n179 gnd.n177 0.00397623
R386 gnd.n70 gnd.n69 0.00391284
R387 gnd.n71 gnd.n70 0.00391159
R388 gnd.n14 gnd.n13 0.00371923
R389 gnd.n11 gnd.n10 0.00294771
R390 gnd.n17 gnd.n16 0.00294771
R391 gnd.n174 gnd.n172 0.00248813
R392 gnd.n258 gnd.n257 0.00245312
R393 gnd.n52 gnd.n51 0.00236777
R394 gnd.n13 gnd.n12 0.00217489
R395 gnd.t111 gnd.n44 0.00192099
R396 gnd.n51 gnd.n50 0.00186816
R397 gnd.n256 gnd.n255 0.00152216
R398 gnd.n169 gnd.n157 0.00152195
R399 gnd.n145 gnd.n137 0.00148887
R400 gnd.n129 gnd.n126 0.00148887
R401 gnd.n215 gnd.n214 0.00138337
R402 gnd.n209 gnd.n208 0.00138109
R403 gnd.n185 gnd.n184 0.00134613
R404 gnd.n179 gnd.n178 0.00134049
R405 gnd.n174 gnd.n173 0.001335
R406 gnd.n50 gnd.n49 0.00124275
R407 gnd.n229 gnd.n228 0.00121065
R408 gnd.n227 gnd.n226 0.001204
R409 gnd.n67 gnd.n66 0.00104118
R410 gnd.n123 gnd.n122 0.00100955
R411 gnd.n68 gnd.n67 0.00100261
R412 gnd.n231 gnd.n230 0.00100079
R413 gnd.n53 gnd.n52 0.00100039
R414 gnd.n203 gnd.n202 0.000522345
R415 gnd.n224 gnd.n223 0.000522345
R416 gnd.n73 gnd.n72 0.00051897
R417 gnd.n216 gnd.n215 0.000501021
R418 gnd.n210 gnd.n209 0.000501021
R419 gnd.n180 gnd.n179 0.000500672
R420 gnd.n186 gnd.n185 0.000500672
R421 buffer_0.a.n6 buffer_0.a.t17 377.647
R422 buffer_0.a.n6 buffer_0.a.t16 376.93
R423 buffer_0.a.n13 buffer_0.a.t4 314.055
R424 buffer_0.a.t0 buffer_0.a.n6 42.2586
R425 buffer_0.a.n7 buffer_0.a.t0 40.2461
R426 buffer_0.a.n1 buffer_0.a.t2 39.5847
R427 buffer_0.a.n11 buffer_0.a.t11 39.5292
R428 buffer_0.a.n9 buffer_0.a.t9 39.5292
R429 buffer_0.a.n8 buffer_0.a.t7 39.5292
R430 buffer_0.a.n7 buffer_0.a.t13 39.5292
R431 buffer_0.a.n2 buffer_0.a.t3 28.5655
R432 buffer_0.a.n2 buffer_0.a.t12 28.5655
R433 buffer_0.a.n3 buffer_0.a.t14 28.5655
R434 buffer_0.a.n3 buffer_0.a.t1 28.5655
R435 buffer_0.a.n4 buffer_0.a.t10 28.5655
R436 buffer_0.a.n4 buffer_0.a.t8 28.5655
R437 buffer_0.a.n13 buffer_0.a.t6 13.2078
R438 buffer_0.a.n0 buffer_0.a.t15 13.2005
R439 buffer_0.a.n0 buffer_0.a.t5 13.2005
R440 buffer_0.a.n5 buffer_0.a.n3 1.62643
R441 buffer_0.a.n10 buffer_0.a.n5 1.438
R442 buffer_0.a.n10 buffer_0.a.n9 1.06207
R443 buffer_0.a.n12 buffer_0.a.n11 1.01015
R444 buffer_0.a.n8 buffer_0.a.n7 0.717388
R445 buffer_0.a.n9 buffer_0.a.n8 0.717388
R446 buffer_0.a buffer_0.a.n0 0.677588
R447 buffer_0.a buffer_0.a.n1 0.45343
R448 buffer_0.a.n5 buffer_0.a.n4 0.157684
R449 buffer_0.a.n0 buffer_0.a.n13 0.119008
R450 buffer_0.a.n11 buffer_0.a.n10 0.0949882
R451 buffer_0.a.n1 buffer_0.a.n12 0.0588333
R452 buffer_0.a.n1 buffer_0.a.n2 0.0587685
R453 sensor_0.b.t8 sensor_0.b.t0 74.8549
R454 sensor_0.b.t6 sensor_0.b.t8 74.8549
R455 sensor_0.b.t14 sensor_0.b.t6 74.8549
R456 sensor_0.b.t10 sensor_0.b.t2 74.8549
R457 sensor_0.b.t4 sensor_0.b.t10 74.8549
R458 sensor_0.b.t12 sensor_0.b.t4 74.8549
R459 sensor_0.b.t24 sensor_0.b.t32 74.8549
R460 sensor_0.b.t31 sensor_0.b.t24 74.8549
R461 sensor_0.b.t23 sensor_0.b.t31 74.8549
R462 sensor_0.b.t34 sensor_0.b.t26 74.8549
R463 sensor_0.b.t21 sensor_0.b.t34 74.8549
R464 sensor_0.b.t29 sensor_0.b.t21 74.8549
R465 sensor_0.b.t27 sensor_0.b.t20 74.8549
R466 sensor_0.b.t28 sensor_0.b.t27 74.8549
R467 sensor_0.b.t35 sensor_0.b.t28 74.8549
R468 sensor_0.b.t22 sensor_0.b.t30 74.8549
R469 sensor_0.b.t33 sensor_0.b.t22 74.8549
R470 sensor_0.b.t25 sensor_0.b.t33 74.8549
R471 sensor_0.b.n7 sensor_0.b.t25 38.3763
R472 sensor_0.b.n11 sensor_0.b.t14 37.3627
R473 sensor_0.b.n10 sensor_0.b.t12 37.3602
R474 sensor_0.b.n9 sensor_0.b.t23 37.3602
R475 sensor_0.b.n8 sensor_0.b.t29 37.3602
R476 sensor_0.b.n7 sensor_0.b.t35 37.3602
R477 sensor_0.b.n12 sensor_0.b.t1 18.2715
R478 sensor_0.b.n3 sensor_0.b.t3 18.1717
R479 sensor_0.b.n14 sensor_0.b.t15 17.427
R480 sensor_0.b.n13 sensor_0.b.t7 17.4116
R481 sensor_0.b.n3 sensor_0.b.t11 17.4101
R482 sensor_0.b.n12 sensor_0.b.t9 17.4101
R483 sensor_0.b.n4 sensor_0.b.t5 17.4058
R484 sensor_0.b.n5 sensor_0.b.t13 17.4056
R485 sensor_0.b.n0 sensor_0.b.t16 14.283
R486 sensor_0.b.n0 sensor_0.b.t18 14.283
R487 sensor_0.b.n1 sensor_0.b.t17 14.283
R488 sensor_0.b.n1 sensor_0.b.t19 14.283
R489 sensor_0.b.n6 sensor_0.b.n5 3.22928
R490 sensor_0.b.n6 sensor_0.b.n2 2.2255
R491 sensor_0.b.n11 sensor_0.b.n10 1.01759
R492 sensor_0.b.n8 sensor_0.b.n7 1.01657
R493 sensor_0.b.n9 sensor_0.b.n8 1.01657
R494 sensor_0.b.n10 sensor_0.b.n9 1.01657
R495 sensor_0.b.n13 sensor_0.b.n12 0.865287
R496 sensor_0.b sensor_0.b.n15 0.851048
R497 sensor_0.b.n14 sensor_0.b.n13 0.777059
R498 sensor_0.b.n5 sensor_0.b.n4 0.718555
R499 sensor_0.b.n4 sensor_0.b.n3 0.710921
R500 sensor_0.b.n2 sensor_0.b.n0 0.49917
R501 sensor_0.b sensor_0.b.n6 0.341125
R502 sensor_0.b.n15 sensor_0.b.n14 0.325292
R503 sensor_0.b.n15 sensor_0.b.n11 0.202053
R504 sensor_0.b.n2 sensor_0.b.n1 0.17167
R505 sensor_0.a.n2 sensor_0.a.t15 64.1667
R506 sensor_0.a.n0 sensor_0.a.t8 63.6292
R507 sensor_0.a.n4 sensor_0.a.t13 63.6292
R508 sensor_0.a.n3 sensor_0.a.t12 63.6292
R509 sensor_0.a.n2 sensor_0.a.t14 63.6292
R510 sensor_0.a.n1 sensor_0.a.t10 63.6275
R511 sensor_0.a.n8 sensor_0.a.t2 18.2715
R512 sensor_0.a.n5 sensor_0.a.t7 18.2714
R513 sensor_0.a.n10 sensor_0.a.t5 17.4132
R514 sensor_0.a.n7 sensor_0.a.t0 17.4132
R515 sensor_0.a.n6 sensor_0.a.t3 17.4116
R516 sensor_0.a.n8 sensor_0.a.t6 17.4101
R517 sensor_0.a.n5 sensor_0.a.t4 17.4101
R518 sensor_0.a.n9 sensor_0.a.t1 17.4057
R519 sensor_0.a.n1 sensor_0.a.t11 14.5343
R520 sensor_0.a.n0 sensor_0.a.t9 14.2976
R521 sensor_0.a sensor_0.a.n11 1.63801
R522 sensor_0.a.n11 sensor_0.a.n7 1.541
R523 sensor_0.a.n11 sensor_0.a.n10 1.541
R524 sensor_0.a.n10 sensor_0.a.n9 0.873387
R525 sensor_0.a.n6 sensor_0.a.n5 0.865287
R526 sensor_0.a.n7 sensor_0.a.n6 0.864262
R527 sensor_0.a.n9 sensor_0.a.n8 0.848309
R528 sensor_0.a.n3 sensor_0.a.n2 0.538
R529 sensor_0.a.n4 sensor_0.a.n3 0.538
R530 sensor_0.a.n0 sensor_0.a.n4 0.488
R531 sensor_0.a.n1 sensor_0.a.n0 0.29354
R532 sensor_0.a sensor_0.a.n1 0.28675
R533 buffer_0.b.n6 buffer_0.b.t17 377.466
R534 buffer_0.b.n6 buffer_0.b.t16 376.93
R535 buffer_0.b.n16 buffer_0.b.t9 313.991
R536 buffer_0.b.t7 buffer_0.b.n6 41.3792
R537 buffer_0.b.n7 buffer_0.b.t7 40.2104
R538 buffer_0.b.n11 buffer_0.b.t13 28.6605
R539 buffer_0.b.n0 buffer_0.b.t15 28.5655
R540 buffer_0.b.n0 buffer_0.b.t12 28.5655
R541 buffer_0.b.n2 buffer_0.b.t8 28.5655
R542 buffer_0.b.n2 buffer_0.b.t6 28.5655
R543 buffer_0.b.n3 buffer_0.b.t4 28.5655
R544 buffer_0.b.n3 buffer_0.b.t2 28.5655
R545 buffer_0.b.n11 buffer_0.b.t11 26.2653
R546 buffer_0.b.n10 buffer_0.b.t14 26.2652
R547 buffer_0.b.n9 buffer_0.b.t1 26.2652
R548 buffer_0.b.n8 buffer_0.b.t3 26.2652
R549 buffer_0.b.n7 buffer_0.b.t5 26.2652
R550 buffer_0.b.n15 buffer_0.b.t0 13.2053
R551 buffer_0.b.n15 buffer_0.b.t10 6.63265
R552 buffer_0.b.n4 buffer_0.b.n2 1.62544
R553 buffer_0.b.n5 buffer_0.b.n4 1.44539
R554 buffer_0.b.n1 buffer_0.b.n10 0.825504
R555 buffer_0.b.n8 buffer_0.b.n7 0.718158
R556 buffer_0.b.n9 buffer_0.b.n8 0.718158
R557 buffer_0.b.n10 buffer_0.b.n9 0.718158
R558 buffer_0.b buffer_0.b.n16 0.594255
R559 buffer_0.b buffer_0.b.n14 0.562809
R560 buffer_0.b.n13 buffer_0.b.n12 0.188
R561 buffer_0.b.n4 buffer_0.b.n3 0.156686
R562 buffer_0.b.n12 buffer_0.b.n1 0.10675
R563 buffer_0.b.n13 buffer_0.b.n5 0.104667
R564 buffer_0.b.n16 buffer_0.b.n15 0.0678366
R565 buffer_0.b.n14 buffer_0.b.n0 0.0624088
R566 buffer_0.b.n1 buffer_0.b.n11 0.0623624
R567 buffer_0.b.n0 buffer_0.b.n13 0.0505
R568 out_buff.n4 out_buff.t3 377.192
R569 out_buff.n1 out_buff.t1 377.175
R570 out_buff.n6 out_buff.t11 317.7
R571 out_buff.n13 out_buff.t6 9.50808
R572 out_buff.n12 out_buff 6.13708
R573 out_buff.n9 out_buff.t5 5.53268
R574 out_buff.n7 out_buff.t0 3.4805
R575 out_buff.n7 out_buff.t7 3.4805
R576 out_buff.n12 out_buff.n11 2.388
R577 out_buff.n5 out_buff.n4 2.02858
R578 out_buff.n2 out_buff.n1 2.00736
R579 out_buff.n3 out_buff.t8 1.90483
R580 out_buff.n3 out_buff.t4 1.90483
R581 out_buff.n0 out_buff.t2 1.90483
R582 out_buff.n0 out_buff.t9 1.90483
R583 out_buff.n6 out_buff.t10 1.78624
R584 out_buff.n8 out_buff.n7 1.58206
R585 out_buff.n13 out_buff.n12 1.11925
R586 out_buff.n10 out_buff.n9 0.80675
R587 out_buff.n9 out_buff.n8 0.770812
R588 out_buff.n11 out_buff.n10 0.722063
R589 out_buff.n10 out_buff.n2 0.182565
R590 out_buff.n9 out_buff.n5 0.182565
R591 out_buff.n11 out_buff 0.06175
R592 out_buff out_buff.n13 0.05675
R593 out_buff.n5 out_buff.n3 0.00195207
R594 out_buff.n2 out_buff.n0 0.00195207
R595 out_buff.n8 out_buff.n6 0.000558569
R596 vd.n61 vd.n43 11483
R597 vd.n56 vd.n43 11371.8
R598 vd.n64 vd.n42 10557.3
R599 vd.n53 vd.n52 10507.9
R600 vd.n45 vd.n42 8128.24
R601 vd.n52 vd.n47 8092.94
R602 vd.n56 vd.n47 6967.06
R603 vd.n61 vd.n45 6931.77
R604 vd.n64 vd.n40 6349.41
R605 vd.n53 vd.n40 6345.88
R606 vd.n18 vd.n15 2142.35
R607 vd.n60 vd.n58 1224.85
R608 vd.n58 vd.n57 1212.99
R609 vd.n22 vd.n16 1164.71
R610 vd.n24 vd.n12 1164.71
R611 vd.n65 vd.n41 1126.12
R612 vd.n50 vd.n39 1120.84
R613 vd.n24 vd.n13 977.648
R614 vd.n22 vd.n15 952.942
R615 vd.n59 vd.n41 867.013
R616 vd.n50 vd.n46 863.247
R617 vd.n57 vd.n46 743.154
R618 vd.n60 vd.n59 739.389
R619 vd.n66 vd.n65 647.907
R620 vd.n66 vd.n39 647.529
R621 vd.t26 vd.t62 331.216
R622 vd.t62 vd.t68 331.216
R623 vd.t68 vd.t66 331.216
R624 vd.t66 vd.t57 331.216
R625 vd.t57 vd.t64 331.216
R626 vd.t64 vd.t61 331.216
R627 vd.t14 vd.t12 331.216
R628 vd.t12 vd.t15 331.216
R629 vd.t15 vd.t6 331.216
R630 vd.t6 vd.t4 331.216
R631 vd.t4 vd.t2 331.216
R632 vd.t2 vd.t29 331.216
R633 vd.n20 vd.n19 228.518
R634 vd.n19 vd.n10 228.518
R635 vd.n48 vd.t14 228.514
R636 vd.t61 vd.n49 210.542
R637 vd.n137 vd.n134 206.306
R638 vd.n105 vd.n104 168.66
R639 vd.t18 vd.n118 156.245
R640 vd.n23 vd.t0 144.606
R641 vd.n100 vd.t38 143.697
R642 vd.n122 vd.t53 143.697
R643 vd.n144 vd.n141 142.306
R644 vd.n18 vd.n17 135.465
R645 vd.n124 vd.n121 126.871
R646 vd.n97 vd.n96 111.421
R647 vd.n25 vd.n10 104.282
R648 vd.n21 vd.n20 101.647
R649 vd.n142 vd.t39 86.6752
R650 vd.n105 vd.n99 85.0829
R651 vd.n135 vd.t22 71.8492
R652 vd.t10 vd.t47 70.1694
R653 vd.t8 vd.t40 70.1694
R654 vd.t42 vd.t59 70.0291
R655 vd.t70 vd.t43 70.0291
R656 vd.n62 vd.t47 68.5376
R657 vd.n100 vd.t33 65.0065
R658 vd.n107 vd.t21 63.9214
R659 vd.n93 vd.t32 63.8352
R660 vd.t40 vd.n42 63.6434
R661 vd.n113 vd.t17 63.6292
R662 vd.n55 vd.t43 63.5148
R663 vd.n137 vd.n131 63.2476
R664 vd.n52 vd.t42 62.9732
R665 vd.n142 vd.t72 60.4447
R666 vd.t39 vd.t36 58.1638
R667 vd.t22 vd.t52 58.1638
R668 vd.n129 vd.t44 42.1974
R669 vd.n132 vd.t51 42.1974
R670 vd.n81 vd.t25 39.5312
R671 vd.n71 vd.t28 39.5292
R672 vd.n49 vd.n48 38.514
R673 vd.n44 vd.t8 37.5327
R674 vd.t59 vd.n51 35.2862
R675 vd.n51 vd.t70 34.7434
R676 vd.n44 vd.t10 32.6372
R677 vd.n26 vd.n25 31.105
R678 vd.t27 vd.n81 28.7267
R679 vd.n71 vd.t31 28.6459
R680 vd.n86 vd.t58 28.5655
R681 vd.n86 vd.t65 28.5655
R682 vd.n82 vd.t27 28.5655
R683 vd.n82 vd.t63 28.5655
R684 vd.n84 vd.t69 28.5655
R685 vd.n84 vd.t67 28.5655
R686 vd.n68 vd.t13 28.5655
R687 vd.n68 vd.t16 28.5655
R688 vd.n70 vd.t3 28.5655
R689 vd.n70 vd.t30 28.5655
R690 vd.n73 vd.t7 28.5655
R691 vd.n73 vd.t5 28.5655
R692 vd.n102 vd.t48 28.5119
R693 vd.n21 vd.n4 27.9188
R694 vd.n115 vd.n110 24.5501
R695 vd.n26 vd.n9 22.401
R696 vd.n34 vd.n33 22.4005
R697 vd.n9 vd.n7 22.4005
R698 vd.n55 vd.n54 21.216
R699 vd.n119 vd.t18 21.0989
R700 vd.t44 vd.t49 19.3883
R701 vd.n35 vd.n4 19.201
R702 vd.n35 vd.n34 19.2005
R703 vd.n135 vd.t50 17.1073
R704 vd.n54 vd.n53 16.7426
R705 vd.n63 vd.t29 16.3842
R706 vd.n63 vd.n62 16.211
R707 vd.n106 vd.t45 14.575
R708 vd.n92 vd.t37 14.5025
R709 vd.n112 vd.t19 14.4041
R710 vd.n94 vd.t34 14.2873
R711 vd.n92 vd.t35 14.2873
R712 vd.n108 vd.t24 14.2873
R713 vd.n106 vd.t23 14.2873
R714 vd.n110 vd.t20 14.2867
R715 vd.n111 vd.t54 14.283
R716 vd.n111 vd.t56 14.283
R717 vd.n54 vd.t26 12.5482
R718 vd.t33 vd.t41 11.4051
R719 vd.n11 vd.n7 10.5605
R720 vd.n33 vd.n6 9.6005
R721 vd.n2 vd.t46 9.5742
R722 vd.n30 vd.t1 9.52337
R723 vd.n115 vd.n114 9.3005
R724 vd.n64 vd.n63 7.64222
R725 vd.n116 vd.n115 4.5005
R726 vd.n75 vd.n67 4.5005
R727 vd.n149 vd.n148 3.79434
R728 vd.n88 vd.n80 3.54402
R729 vd.n79 vd.n78 3.47391
R730 vd.n122 vd.t55 3.42187
R731 vd vd.n38 2.438
R732 vd.n11 vd.n6 2.2405
R733 vd.n80 vd.t60 1.90483
R734 vd.n80 vd.t71 1.90483
R735 vd.n78 vd.t11 1.90483
R736 vd.n78 vd.t9 1.90483
R737 vd vd.n116 1.83279
R738 vd.n91 vd 1.73266
R739 vd.n85 vd.n83 1.56925
R740 vd.n74 vd.n72 1.5417
R741 vd.n87 vd.n85 1.44593
R742 vd.n75 vd.n74 1.38331
R743 vd.n147 vd.n94 0.881455
R744 vd.n148 vd.n147 0.834744
R745 vd.n112 vd.n111 0.721906
R746 vd.n83 vd.n81 0.686006
R747 vd.n113 vd.n112 0.608294
R748 vd.n126 vd.n108 0.59946
R749 vd.n146 vd.n145 0.5755
R750 vd.n89 vd.n79 0.497524
R751 vd.n145 vd.n138 0.488
R752 vd.n126 vd.n125 0.463
R753 vd.n89 vd.n88 0.4255
R754 vd.n88 vd.n87 0.424134
R755 vd.n148 vd.n91 0.328325
R756 vd.n79 vd.n77 0.313286
R757 vd.n125 vd 0.2755
R758 vd.n138 vd.n126 0.238
R759 vd.n150 vd.n149 0.2005
R760 vd.n85 vd.n84 0.157684
R761 vd.n74 vd.n73 0.156686
R762 vd.n28 vd.n27 0.146341
R763 vd.n28 vd.n3 0.146333
R764 vd.n107 vd.n106 0.134875
R765 vd.n108 vd.n107 0.134875
R766 vd.n22 vd.n21 0.130052
R767 vd.n23 vd.n22 0.130052
R768 vd.n38 vd.n3 0.1255
R769 vd.n150 vd 0.1255
R770 vd.n110 vd.n109 0.122252
R771 vd.n114 vd.n113 0.116172
R772 vd.n94 vd.n93 0.115679
R773 vd.n93 vd.n92 0.115679
R774 vd.n25 vd.n24 0.107375
R775 vd.n24 vd.n23 0.107375
R776 vd.n91 vd 0.100725
R777 vd.n150 vd.n2 0.0822638
R778 vd.n72 vd.n71 0.0791768
R779 vd.n0 vd.t73 0.0686501
R780 vd.n1 vd.n0 0.06865
R781 vd.n72 vd.n70 0.0493677
R782 vd.n76 vd.n75 0.0489375
R783 vd.n83 vd.n82 0.0461626
R784 vd.n32 vd.n5 0.0456031
R785 vd.n29 vd.n8 0.0456031
R786 vd.n27 vd.n8 0.0456031
R787 vd.n37 vd.n36 0.0391598
R788 vd.n36 vd.n5 0.0391598
R789 vd.n149 vd 0.0372647
R790 vd.n20 vd.n15 0.0349892
R791 vd.n15 vd.t0 0.0349892
R792 vd.n13 vd.n10 0.0349892
R793 vd vd.n90 0.0347717
R794 vd.n17 vd.n13 0.0333079
R795 vd.n99 vd.n98 0.0307238
R796 vd.n98 vd.n97 0.0302348
R797 vd.n30 vd.n29 0.0217629
R798 vd.n69 vd.n68 0.0200317
R799 vd.n32 vd.n31 0.0198299
R800 vd.n77 vd.n67 0.01975
R801 vd.n116 vd.n109 0.0176875
R802 vd.n121 vd.n120 0.0175052
R803 vd.n120 vd.n119 0.0175052
R804 vd.n141 vd.n140 0.0150968
R805 vd.n140 vd.n139 0.0150968
R806 vd.n87 vd.n86 0.0148061
R807 vd.n69 vd.n67 0.0141783
R808 vd vd.n150 0.013
R809 vd.n14 vd.n12 0.0125538
R810 vd.n104 vd.n103 0.0122827
R811 vd.n103 vd.n102 0.0122827
R812 vd.n12 vd.n11 0.0120596
R813 vd.n114 vd.n109 0.009875
R814 vd.n134 vd.n133 0.00973799
R815 vd.n133 vd.n132 0.00973799
R816 vd.n2 vd.n1 0.00846782
R817 vd.n76 vd.n69 0.0083125
R818 vd.n147 vd.n146 0.00675
R819 vd.n19 vd.n18 0.00627981
R820 vd.n31 vd.n30 0.00501031
R821 vd.n47 vd.n46 0.00431884
R822 vd.n51 vd.n47 0.00431884
R823 vd.n59 vd.n45 0.00425193
R824 vd.n45 vd.n44 0.00425193
R825 vd.n144 vd.n143 0.00391284
R826 vd.n143 vd.n142 0.00391284
R827 vd.n137 vd.n136 0.00391284
R828 vd.n136 vd.n135 0.00391284
R829 vd.n124 vd.n123 0.00391284
R830 vd.n123 vd.n122 0.00391284
R831 vd.n105 vd.n101 0.00391284
R832 vd.n101 vd.n100 0.00391284
R833 vd.n65 vd.n64 0.00389051
R834 vd.n53 vd.n39 0.00389051
R835 vd.n118 vd.n117 0.00347027
R836 vd.n96 vd.n95 0.00347027
R837 vd.n17 vd.t0 0.00318081
R838 vd.n131 vd.n130 0.00275116
R839 vd.n130 vd.n129 0.00275116
R840 vd.n61 vd.n60 0.0021559
R841 vd.n62 vd.n61 0.0021559
R842 vd.n57 vd.n56 0.00213065
R843 vd.n56 vd.n55 0.00213065
R844 vd.n90 vd.n66 0.00200289
R845 vd.n16 vd.n14 0.0018171
R846 vd.n42 vd.n41 0.00181202
R847 vd.n52 vd.n50 0.00181202
R848 vd.n58 vd.n43 0.0017783
R849 vd.n49 vd.n43 0.0017783
R850 vd.n129 vd.n128 0.00162558
R851 vd.n128 vd.n127 0.00162558
R852 vd.n16 vd.n6 0.00131751
R853 vd.n31 vd.n6 0.00131744
R854 vd.n36 vd.n35 0.00119114
R855 vd.n37 vd.n4 0.00101609
R856 vd.n77 vd.n76 0.00100557
R857 vd.n90 vd.n89 0.00100109
R858 vd.n23 vd.n14 0.00100038
R859 vd.n27 vd.n26 0.00100009
R860 vd.n66 vd.n40 0.000827345
R861 vd.n48 vd.n40 0.000827345
R862 vd.n9 vd.n8 0.000659706
R863 vd.n33 vd.n32 0.000659706
R864 vd.n34 vd.n5 0.000543686
R865 vd.n29 vd.n7 0.000543686
R866 vd.n145 vd.n144 0.000532663
R867 vd.n138 vd.n137 0.000532663
R868 vd.n125 vd.n124 0.000532663
R869 vd.n146 vd.n105 0.000532663
R870 vd.n38 vd.n37 0.000507883
R871 vd.n5 vd.n3 0.000507883
R872 vd.n29 vd.n28 0.000507883
R873 vd.n0 vd.t75 0.000500086
R874 vd.n1 vd.t74 0.000500086
R875 vpwr.t17 vpwr.t20 790.188
R876 vpwr.t4 vpwr.t0 648.131
R877 vpwr.t26 vpwr.t6 583.023
R878 vpwr.n77 vpwr 548.548
R879 vpwr.n56 vpwr.t7 514.011
R880 vpwr.t14 vpwr.t4 485.358
R881 vpwr.t16 vpwr.t28 414.33
R882 vpwr.n14 vpwr.t25 413.315
R883 vpwr.n32 vpwr.t21 375.277
R884 vpwr.n7 vpwr.t22 344.005
R885 vpwr.t2 vpwr.t23 319.627
R886 vpwr.n50 vpwr.n39 311.957
R887 vpwr.n72 vpwr.n31 311.894
R888 vpwr.n59 vpwr.n58 309.18
R889 vpwr.t6 vpwr.t19 292.991
R890 vpwr.t8 vpwr.t16 292.991
R891 vpwr.n43 vpwr.n40 292.5
R892 vpwr.n45 vpwr.n44 292.5
R893 vpwr.t0 vpwr.t10 287.072
R894 vpwr.t28 vpwr.t26 287.072
R895 vpwr.t20 vpwr.t8 272.274
R896 vpwr.t19 vpwr.t9 254.518
R897 vpwr.t23 vpwr.t14 248.599
R898 vpwr.t9 vpwr.t2 248.599
R899 vpwr.t12 vpwr.t17 244.306
R900 vpwr.n6 vpwr.t31 187.321
R901 vpwr vpwr.t12 186.556
R902 vpwr.n44 vpwr.n43 182.929
R903 vpwr.n7 vpwr.n5 152
R904 vpwr.n42 vpwr.n41 148.689
R905 vpwr.n14 vpwr.t30 126.127
R906 vpwr.n39 vpwr.t3 119.608
R907 vpwr.n58 vpwr.t29 93.81
R908 vpwr.n6 vpwr.n1 73.2067
R909 vpwr.n43 vpwr.t15 68.0124
R910 vpwr.n58 vpwr.t27 63.3219
R911 vpwr.n39 vpwr.t24 63.3219
R912 vpwr.n41 vpwr.t1 61.9158
R913 vpwr.n31 vpwr.t18 41.5552
R914 vpwr.n31 vpwr.t13 41.5552
R915 vpwr.n71 vpwr.n70 34.6358
R916 vpwr.n64 vpwr.n34 34.6358
R917 vpwr.n65 vpwr.n64 34.6358
R918 vpwr.n66 vpwr.n65 34.6358
R919 vpwr.n60 vpwr.n57 34.6358
R920 vpwr.n51 vpwr.n37 34.6358
R921 vpwr.n55 vpwr.n37 34.6358
R922 vpwr.n66 vpwr.n32 32.377
R923 vpwr.n56 vpwr.n55 32.0005
R924 vpwr.n41 vpwr.t11 30.239
R925 vpwr.n50 vpwr.n49 30.1181
R926 vpwr.n44 vpwr.t5 29.316
R927 vpwr.n72 vpwr.n71 22.9652
R928 vpwr.n51 vpwr.n50 20.3299
R929 vpwr.n70 vpwr.n32 18.0711
R930 vpwr vpwr.n4 14.0185
R931 vpwr.n45 vpwr.n42 13.9946
R932 vpwr.n49 vpwr.n40 12.8758
R933 vpwr.n57 vpwr.n56 9.41227
R934 vpwr.n11 vpwr.n10 9.3005
R935 vpwr.n8 vpwr.n2 9.3005
R936 vpwr.n8 vpwr.n7 9.3005
R937 vpwr.n7 vpwr.n6 9.15991
R938 vpwr.n15 vpwr.n14 7.02651
R939 vpwr.n59 vpwr.n34 6.02403
R940 vpwr.n46 vpwr.n45 5.00414
R941 vpwr.n4 vpwr 4.7293
R942 vpwr.n9 vpwr.n0 4.6505
R943 vpwr.n18 vpwr.n17 4.6505
R944 vpwr.n47 vpwr.n46 4.6505
R945 vpwr.n49 vpwr.n48 4.6505
R946 vpwr.n50 vpwr.n38 4.6505
R947 vpwr.n52 vpwr.n51 4.6505
R948 vpwr.n53 vpwr.n37 4.6505
R949 vpwr.n55 vpwr.n54 4.6505
R950 vpwr.n56 vpwr.n36 4.6505
R951 vpwr.n57 vpwr.n35 4.6505
R952 vpwr.n61 vpwr.n60 4.6505
R953 vpwr.n62 vpwr.n34 4.6505
R954 vpwr.n64 vpwr.n63 4.6505
R955 vpwr.n65 vpwr.n33 4.6505
R956 vpwr.n67 vpwr.n66 4.6505
R957 vpwr.n68 vpwr.n32 4.6505
R958 vpwr.n70 vpwr.n69 4.6505
R959 vpwr.n71 vpwr.n30 4.6505
R960 vpwr.n4 vpwr 4.53383
R961 vpwr.n46 vpwr.n40 4.07323
R962 vpwr.n73 vpwr.n72 3.93272
R963 vpwr.n60 vpwr.n59 3.76521
R964 vpwr.n5 vpwr 3.11401
R965 vpwr.n17 vpwr.n15 3.0725
R966 vpwr.n28 vpwr 2.92878
R967 vpwr.n27 vpwr.n26 2.91783
R968 vpwr.n12 vpwr 2.36657
R969 vpwr.n5 vpwr.n1 1.55726
R970 vpwr.n10 vpwr.n9 1.55726
R971 vpwr.n8 vpwr.n1 1.38428
R972 vpwr.n9 vpwr.n8 1.38428
R973 vpwr.n10 vpwr 1.38428
R974 vpwr.n17 vpwr.n16 1.2805
R975 vpwr.n77 vpwr.n76 0.711611
R976 vpwr.n12 vpwr 0.580857
R977 vpwr.n29 vpwr.n28 0.5255
R978 vpwr.n75 vpwr 0.223
R979 vpwr.n3 vpwr 0.196446
R980 vpwr.n20 vpwr 0.171696
R981 vpwr.n47 vpwr.n42 0.144332
R982 vpwr.n73 vpwr.n30 0.138831
R983 vpwr.n48 vpwr.n47 0.120292
R984 vpwr.n48 vpwr.n38 0.120292
R985 vpwr.n52 vpwr.n38 0.120292
R986 vpwr.n53 vpwr.n52 0.120292
R987 vpwr.n54 vpwr.n53 0.120292
R988 vpwr.n54 vpwr.n36 0.120292
R989 vpwr.n36 vpwr.n35 0.120292
R990 vpwr.n61 vpwr.n35 0.120292
R991 vpwr.n62 vpwr.n61 0.120292
R992 vpwr.n63 vpwr.n62 0.120292
R993 vpwr.n63 vpwr.n33 0.120292
R994 vpwr.n67 vpwr.n33 0.120292
R995 vpwr.n68 vpwr.n67 0.120292
R996 vpwr.n69 vpwr.n68 0.120292
R997 vpwr.n69 vpwr.n30 0.120292
R998 vpwr.n74 vpwr.n73 0.107496
R999 vpwr.n20 vpwr.n19 0.0901739
R1000 vpwr vpwr.n83 0.0634013
R1001 vpwr.n27 vpwr 0.063
R1002 vpwr.n21 vpwr.n20 0.0500874
R1003 vpwr.n13 vpwr.n12 0.0466957
R1004 vpwr.n24 vpwr.n23 0.0435328
R1005 vpwr.n83 vpwr.n29 0.039096
R1006 vpwr.n18 vpwr.n13 0.0331087
R1007 vpwr.n83 vpwr.n82 0.0287348
R1008 vpwr.n3 vpwr.n2 0.02675
R1009 vpwr vpwr.n11 0.0255
R1010 vpwr.n22 vpwr.n21 0.0213989
R1011 vpwr.n78 vpwr.n75 0.0207266
R1012 vpwr.n26 vpwr.n25 0.018111
R1013 vpwr.n74 vpwr 0.0174271
R1014 vpwr vpwr.n74 0.01675
R1015 vpwr.n19 vpwr.n18 0.014087
R1016 vpwr.n24 vpwr.n22 0.0127951
R1017 vpwr.n11 vpwr.n0 0.01175
R1018 vpwr.n2 vpwr.n0 0.0105
R1019 vpwr.n81 vpwr.n80 0.009875
R1020 vpwr vpwr.n3 0.00725676
R1021 vpwr.n23 vpwr 0.00459836
R1022 vpwr.n79 vpwr.n78 0.00412592
R1023 vpwr.n80 vpwr.n79 0.003625
R1024 vpwr.n82 vpwr.n81 0.00196888
R1025 vpwr.n26 vpwr.n24 0.0016109
R1026 vpwr.n78 vpwr.n77 0.00154933
R1027 vpwr.n28 vpwr.n27 0.000500433
R1028 vtd.n7 vtd.t29 64.6821
R1029 vtd.n8 vtd.t27 64.3461
R1030 vtd.n4 vtd.t24 63.6317
R1031 vtd.n9 vtd.t26 63.6292
R1032 vtd.n8 vtd.t28 63.6292
R1033 vtd.n17 vtd.t14 63.6292
R1034 vtd.n2 vtd.t16 63.6292
R1035 vtd.n18 vtd.t22 63.6292
R1036 vtd.n1 vtd.t8 63.6292
R1037 vtd.n19 vtd.t12 63.6292
R1038 vtd.n0 vtd.t18 63.6292
R1039 vtd.n6 vtd.t20 63.6292
R1040 vtd.n3 vtd.t10 63.6275
R1041 vtd.n13 vtd.t4 18.2948
R1042 vtd.n10 vtd.t1 18.1899
R1043 vtd.n10 vtd.t5 17.4187
R1044 vtd.n13 vtd.t0 17.4177
R1045 vtd.n11 vtd.t2 17.4156
R1046 vtd.n14 vtd.t7 17.4136
R1047 vtd.n12 vtd.t6 17.4125
R1048 vtd.n15 vtd.t3 17.4115
R1049 vtd.n3 vtd.t11 14.3559
R1050 vtd.n17 vtd.t15 14.3555
R1051 vtd.n2 vtd.t23 14.283
R1052 vtd.n2 vtd.t17 14.283
R1053 vtd.n1 vtd.t13 14.283
R1054 vtd.n1 vtd.t9 14.283
R1055 vtd.n0 vtd.t21 14.283
R1056 vtd.n0 vtd.t19 14.283
R1057 vtd.n7 vtd.t25 13.7801
R1058 vtd.n16 vtd.n15 2.14635
R1059 vtd.n3 vtd.n16 1.54335
R1060 vtd vtd.n20 1.22372
R1061 vtd.n16 vtd.n12 1.09526
R1062 vtd.n20 vtd.n3 0.981002
R1063 vtd.n15 vtd.n14 0.8755
R1064 vtd.n14 vtd.n13 0.8755
R1065 vtd.n5 vtd.n7 0.832184
R1066 vtd.n11 vtd.n10 0.769433
R1067 vtd.n12 vtd.n11 0.769356
R1068 vtd.n9 vtd.n8 0.717388
R1069 vtd.n4 vtd.n9 0.708453
R1070 vtd.n20 vtd.n5 0.438348
R1071 vtd.n3 vtd.n6 0.140567
R1072 vtd.n18 vtd.n2 0.140142
R1073 vtd.n19 vtd.n1 0.140142
R1074 vtd.n6 vtd.n0 0.140142
R1075 vtd.n0 vtd.n19 0.134875
R1076 vtd.n1 vtd.n18 0.134875
R1077 vtd.n2 vtd.n17 0.134875
R1078 vtd.n5 vtd.n4 0.114328
R1079 buffer_0.d.n9 buffer_0.d.t4 377.216
R1080 buffer_0.d.n8 buffer_0.d.t2 377.163
R1081 buffer_0.d.n2 buffer_0.d.t12 134.298
R1082 buffer_0.d.n4 buffer_0.d.t7 133.787
R1083 buffer_0.d.n3 buffer_0.d.t9 133.761
R1084 buffer_0.d.n2 buffer_0.d.t13 133.761
R1085 buffer_0.d.n1 buffer_0.d.t6 5.55126
R1086 buffer_0.d.n6 buffer_0.d.t10 3.4805
R1087 buffer_0.d.n6 buffer_0.d.t8 3.4805
R1088 buffer_0.d buffer_0.d.n7 3.10062
R1089 buffer_0.d.n1 buffer_0.d.n9 2.02586
R1090 buffer_0.d.n0 buffer_0.d.n8 1.99422
R1091 buffer_0.d.n5 buffer_0.d.t11 1.91167
R1092 buffer_0.d.n0 buffer_0.d.t1 1.9057
R1093 buffer_0.d.n1 buffer_0.d.t0 1.90483
R1094 buffer_0.d.n1 buffer_0.d.t5 1.90483
R1095 buffer_0.d.n0 buffer_0.d.t3 1.42659
R1096 buffer_0.d buffer_0.d.n0 0.77675
R1097 buffer_0.d.n0 buffer_0.d.n1 0.648539
R1098 buffer_0.d.n3 buffer_0.d.n2 0.538
R1099 buffer_0.d.n4 buffer_0.d.n3 0.394346
R1100 buffer_0.d.n7 buffer_0.d.n6 0.151643
R1101 buffer_0.d.n5 buffer_0.d.n4 0.0558728
R1102 buffer_0.d.n7 buffer_0.d.n5 0.0333947
R1103 ib.n0 ib.t5 38.0465
R1104 ib.n0 ib.t3 37.3602
R1105 ib.n4 ib.t0 18.7496
R1106 ib.n4 ib.t2 17.4934
R1107 ib.n1 ib.t4 17.4005
R1108 ib.n1 ib.t1 17.4005
R1109 ib.n9 ib.n8 5.70556
R1110 ib.n3 ib.n2 1.98477
R1111 ib.n8 ib.n0 0.247263
R1112 ib.n10 ib 0.129406
R1113 ib.n9 ib 0.1205
R1114 ib.n5 ib.n4 0.102062
R1115 ib ib.n10 0.0605
R1116 ib.n8 ib.n7 0.059593
R1117 ib.n7 ib.n6 0.0239375
R1118 ib.n6 ib.n3 0.0166802
R1119 ib.n6 ib.n5 0.003625
R1120 ib.n3 ib.n1 0.00322924
R1121 ib.n10 ib.n9 0.00114405
R1122 vts.n23 vts.n18 761.601
R1123 vts.n24 vts.n23 641.883
R1124 vts.t18 vts.t5 333.303
R1125 vts.n35 vts.t25 325.759
R1126 vts.n17 vts.t22 262.014
R1127 vts.n26 vts.t18 237.054
R1128 vts.t5 vts.t2 229.925
R1129 vts.t15 vts.t0 229.925
R1130 vts.t13 vts.t11 229.925
R1131 vts.t11 vts.t9 229.925
R1132 vts.t9 vts.t7 229.925
R1133 vts.n21 vts.t15 130.113
R1134 vts.n21 vts.t13 99.8129
R1135 vts.n11 vts.t17 63.6292
R1136 vts.n4 vts.t21 63.6292
R1137 vts.n31 vts.t4 16.8006
R1138 vts.n5 vts.t23 14.4639
R1139 vts.n10 vts.t20 14.4362
R1140 vts.n12 vts.t19 14.4313
R1141 vts.n4 vts.t24 14.3697
R1142 vts.n0 vts.t6 14.283
R1143 vts.n0 vts.t3 14.283
R1144 vts.n1 vts.t1 14.283
R1145 vts.n1 vts.t16 14.283
R1146 vts.n2 vts.t14 14.283
R1147 vts.n2 vts.t12 14.283
R1148 vts.n3 vts.t10 14.283
R1149 vts.n3 vts.t8 14.283
R1150 vts.n36 vts 3.48645
R1151 vts.n36 vts.n35 1.21925
R1152 vts vts.n34 0.8255
R1153 vts.n9 vts.n8 0.6455
R1154 vts.n8 vts.n7 0.6455
R1155 vts.n7 vts.n6 0.6455
R1156 vts.n6 vts.n5 0.450361
R1157 vts.n10 vts.n9 0.440551
R1158 vts vts.n36 0.26925
R1159 vts.n30 vts.n12 0.0947919
R1160 vts.n5 vts.n4 0.0741592
R1161 vts.n11 vts.n10 0.0682354
R1162 vts.n12 vts.n11 0.0634447
R1163 vts.n35 vts 0.058
R1164 vts.n34 vts.n33 0.05093
R1165 vts.n25 vts.n24 0.0426316
R1166 vts.n26 vts.n25 0.0426316
R1167 vts.n16 vts.n15 0.0175052
R1168 vts.n26 vts.n16 0.0175052
R1169 vts.n9 vts.n0 0.0129196
R1170 vts.n8 vts.n1 0.0129196
R1171 vts.n7 vts.n2 0.0129196
R1172 vts.n6 vts.n3 0.0129196
R1173 vts.n27 vts.n14 0.011183
R1174 vts.n14 vts.n13 0.0106833
R1175 vts.n28 vts.n27 0.0075124
R1176 vts.n29 vts.n28 0.00701261
R1177 vts.n18 vts.n17 0.00559165
R1178 vts.n23 vts.n22 0.00192573
R1179 vts.n22 vts.n21 0.00192573
R1180 vts.n20 vts.n19 0.00192573
R1181 vts.n21 vts.n20 0.00192573
R1182 vts.n33 vts.n32 0.00151802
R1183 vts.n32 vts.n30 0.00150795
R1184 vts.n27 vts.n26 0.00100013
R1185 vts.n30 vts.n29 0.00100001
R1186 vts.n32 vts.n31 0.001
R1187 out_sigma.n1 out_sigma.t2 394.808
R1188 out_sigma.n0 out_sigma.t1 250.941
R1189 out_sigma out_sigma.t0 144.601
R1190 out_sigma out_sigma.n1 9.0826
R1191 out_sigma out_sigma.n0 4.7225
R1192 out_sigma.n2 out_sigma 4.48083
R1193 out_sigma.n0 out_sigma 3.35288
R1194 out_sigma.n2 out_sigma 3.2272
R1195 out_sigma.n1 out_sigma 0.727062
R1196 out_sigma out_sigma.n2 0.13175
R1197 clk.n0 clk.t0 294.557
R1198 clk.n0 clk.t1 211.01
R1199 clk.n2 clk.n0 8.28655
R1200 clk.n3 clk 7.73487
R1201 clk.n3 clk.n2 1.82961
R1202 clk.n1 clk 0.981259
R1203 clk.n2 clk.n1 0.848973
R1204 clk clk.n5 0.385917
R1205 clk.n5 clk.n4 0.03175
R1206 clk.n4 clk.n3 0.00111796
R1207 out.n2 out.t0 8.97158
R1208 out.n2 out.n1 2.56714
R1209 out.n0 out.t2 0.506271
R1210 out.n1 out.n0 0.504061
R1211 out out.n2 0.240344
R1212 out.n0 out.t1 0.0277714
R1213 out.n1 out.t3 0.00303875
C0 sigma-delta_0.x1.Q vd 0.0969f
C1 a_14791_2515# out_sigma 0.00128f
C2 vd a_6126_29386# 0.0189f
C3 vpwr a_16445_2515# 0.2f
C4 ib buffer_0.c 0.185f
C5 out a_16688_5320# 0.00185f
C6 sensor_0.c vts 0.166f
C7 a_16356_5320# out 0.00195f
C8 a_16024_5320# a_15546_5320# 0.144f
C9 buffer_0.a buffer_0.b 0.239f
C10 out_buff out 0.00558f
C11 out a_15214_5320# 0.00184f
C12 sigma-delta_0.x1.Q a_15712_3988# 0.414f
C13 a_16688_5320# a_16854_3988# 0.00473f
C14 a_16445_2515# a_16522_3988# 1.4e-19
C15 sensor_0.a vts 0.543f
C16 a_14791_2515# vd 1.08e-19
C17 sigma-delta_0.x1.Q a_17020_5320# 0.00839f
C18 out_buff clk 0.865f
C19 buffer_0.a buffer_0.c 0.199f
C20 sigma-delta_0.x1.Q a_15141_2515# 8.11e-19
C21 a_16060_2515# sigma-delta_0.x1.Q 6.05e-19
C22 a_14625_2515# sigma-delta_0.x1.Q 9.54e-19
C23 vd a_16190_3988# 0.00388f
C24 a_15546_5320# out 0.00187f
C25 out_buff a_15048_3988# 0.00138f
C26 a_15706_2515# a_16445_2515# 7.05e-19
C27 a_15048_3988# a_15214_5320# 0.00473f
C28 out_buff a_14550_5320# 0.0535f
C29 a_15046_2515# clk 3.09e-19
C30 out_buff sigma-delta_0.x1.D 1.65e-19
C31 a_14791_2515# a_15712_3988# 4.13e-19
C32 vpwr sigma-delta_0.x1.Q 0.186f
C33 clk a_15815_2515# 1.1e-20
C34 out_sigma vd 1.06f
C35 a_15237_2515# sigma-delta_0.x1.Q 1.45e-19
C36 out_buff vts 0.103f
C37 buffer_0.d out 5.5e-19
C38 a_14791_2515# a_15141_2515# 0.23f
C39 a_16190_3988# a_15712_3988# 0.357f
C40 a_14625_2515# a_14791_2515# 0.906f
C41 a_15046_2515# sigma-delta_0.x1.D 0.164f
C42 sigma-delta_0.x1.Q a_16522_3988# 5e-20
C43 a_15249_2881# a_15359_2757# 0.0977f
C44 buffer_0.d clk 0.109f
C45 sigma-delta_0.x1.D a_15815_2515# 2.42e-20
C46 sigma-delta_0.x1.Q a_15403_2515# 9.75e-20
C47 a_15359_2757# clk 1.78e-19
C48 out_sigma a_15712_3988# 0.16f
C49 vpwr a_14791_2515# 0.607f
C50 sigma-delta_0.x1.Q a_15706_2515# 0.00593f
C51 a_15237_2515# a_14791_2515# 2.28e-19
C52 a_15868_2881# a_15359_2757# 2.6e-19
C53 out_sigma buffer_0.b 0.0176f
C54 sigma-delta_0.x1.Q a_15380_3988# 1.43e-21
C55 out_sigma a_15141_2515# 7.05e-19
C56 vpwr a_16190_3988# 0.00384f
C57 a_14625_2515# out_sigma 0.00261f
C58 a_16024_5320# out 0.00189f
C59 sigma-delta_0.x1.D a_15359_2757# 6.24e-19
C60 vd a_15712_3988# 0.75f
C61 sensor_0.d vd 0.282f
C62 vd buffer_0.b 6.27f
C63 vd a_17020_5320# 0.201f
C64 buffer_0.d vts 0.832f
C65 a_15048_3988# a_14716_3988# 0.296f
C66 out_buff ib 0.112f
C67 a_16522_3988# a_16190_3988# 0.312f
C68 vpwr out_sigma 2.26f
C69 a_14625_2515# vd 1.72e-20
C70 a_14716_3988# a_14550_5320# 0.00458f
C71 a_14791_2515# a_15706_2515# 0.125f
C72 vd a_14882_5320# 0.061f
C73 sigma-delta_0.x1.D a_14716_3988# 2.07e-19
C74 vd buffer_0.c 0.00573f
C75 vpwr vd 0.00726f
C76 a_17020_5320# a_15712_3988# 0.00974f
C77 buffer_0.a out_buff 0.0961f
C78 a_15712_3988# a_15141_2515# 2.02e-20
C79 sigma-delta_0.x1.Q a_16688_5320# 0.0032f
C80 sensor_0.b vts 1f
C81 a_14625_2515# a_15712_3988# 1.78e-19
C82 out_sigma a_15706_2515# 6.85e-19
C83 out_sigma a_15380_3988# 0.0148f
C84 vd a_16522_3988# 0.00558f
C85 out a_14550_5320# 0.00197f
C86 a_14625_2515# a_15141_2515# 0.115f
C87 buffer_0.b buffer_0.c 0.16f
C88 buffer_0.d ib 0.766f
C89 vpwr a_15712_3988# 0.0132f
C90 a_15249_2881# sigma-delta_0.x1.D 5.56e-20
C91 a_15046_2515# sigma-delta_0.x1.Q 7.58e-20
C92 clk a_15881_2489# 2.68e-20
C93 vd a_15706_2515# 3.52e-19
C94 vd a_15380_3988# 0.00209f
C95 sigma-delta_0.x1.D a_16854_3988# 2.69e-19
C96 sigma-delta_0.x1.D clk 0.00993f
C97 vpwr a_15141_2515# 0.363f
C98 vpwr a_16060_2515# 0.00312f
C99 sigma-delta_0.x1.Q a_15815_2515# 1.47e-19
C100 a_15237_2515# a_15141_2515# 0.0138f
C101 vpwr a_14625_2515# 0.772f
C102 sensor_0.c vd 0.804f
C103 a_15868_2881# sigma-delta_0.x1.D 2.11e-20
C104 a_15237_2515# a_14625_2515# 0.00134f
C105 out_buff a_14791_2515# 8.29e-20
C106 a_16522_3988# a_15712_3988# 0.0502f
C107 sigma-delta_0.x1.D a_15048_3988# 2.56e-20
C108 buffer_0.a buffer_0.d 1.27f
C109 a_16356_5320# a_16190_3988# 0.00536f
C110 sigma-delta_0.x1.D a_15881_2489# 0.004f
C111 out_buff a_16190_3988# 9.87e-22
C112 sensor_0.a vd 2.92f
C113 a_15403_2515# a_15141_2515# 0.00171f
C114 a_15706_2515# a_15712_3988# 0.0011f
C115 a_15237_2515# vpwr 0.00292f
C116 a_15712_3988# a_15380_3988# 0.298f
C117 a_15046_2515# a_14791_2515# 0.0642f
C118 a_15359_2757# sigma-delta_0.x1.Q 0.00111f
C119 a_14791_2515# a_15815_2515# 2.36e-20
C120 a_15706_2515# a_15141_2515# 7.99e-20
C121 sensor_0.d sensor_0.c 0.492f
C122 a_15380_3988# a_15141_2515# 1.22e-19
C123 out_buff out_sigma 2.45f
C124 a_14625_2515# a_15706_2515# 0.102f
C125 vpwr a_16522_3988# 0.00266f
C126 vpwr a_15403_2515# 0.00407f
C127 vd a_16688_5320# 0.0633f
C128 sensor_0.d sensor_0.a 0.588f
C129 vd a_16356_5320# 0.0637f
C130 vpwr a_15706_2515# 0.524f
C131 out_buff vd 5.19f
C132 vpwr a_15380_3988# 0.00397f
C133 a_14791_2515# a_15359_2757# 0.186f
C134 vd a_15214_5320# 0.0598f
C135 a_16445_2515# a_15881_2489# 0.107f
C136 sigma-delta_0.x1.D a_16445_2515# 0.00209f
C137 buffer_0.a out 0.00222f
C138 a_16688_5320# a_15712_3988# 0.00557f
C139 vd a_15546_5320# 0.0619f
C140 a_16356_5320# a_15712_3988# 0.00631f
C141 a_17020_5320# a_16688_5320# 0.299f
C142 buffer_0.d out_sigma 0.00232f
C143 out_buff a_15712_3988# 0.00915f
C144 a_15359_2757# out_sigma 3.73e-19
C145 out_buff buffer_0.b 2.01f
C146 a_15249_2881# sigma-delta_0.x1.Q 3.66e-19
C147 ib vts 1.08f
C148 a_6126_29386# out 0.0171f
C149 sigma-delta_0.x1.Q a_16854_3988# 0.414f
C150 out_buff a_14625_2515# 4.76e-19
C151 a_16024_5320# a_16190_3988# 0.00473f
C152 out_buff a_14882_5320# 0.0014f
C153 buffer_0.d vd 4.12f
C154 a_15868_2881# sigma-delta_0.x1.Q 4.53e-20
C155 out_buff buffer_0.c 0.0405f
C156 a_15546_5320# a_15712_3988# 0.00466f
C157 a_15214_5320# a_14882_5320# 0.303f
C158 out_sigma a_14716_3988# 0.0146f
C159 a_15815_2515# a_15712_3988# 1.36e-20
C160 a_15046_2515# a_15141_2515# 0.0498f
C161 sigma-delta_0.x1.Q a_15881_2489# 0.142f
C162 out_buff vpwr 0.0121f
C163 a_15046_2515# a_14625_2515# 0.0931f
C164 sigma-delta_0.x1.D sigma-delta_0.x1.Q 0.0675f
C165 buffer_0.a vts 0.253f
C166 sensor_0.c sensor_0.a 0.997f
C167 a_15249_2881# a_14791_2515# 0.0346f
C168 a_14625_2515# a_15815_2515# 2.56e-19
C169 a_16688_5320# a_16522_3988# 0.00482f
C170 vd a_14716_3988# 0.0021f
C171 a_16356_5320# a_16522_3988# 0.00509f
C172 a_14791_2515# clk 0.00241f
C173 buffer_0.d buffer_0.b 0.0351f
C174 vpwr a_15046_2515# 0.0861f
C175 a_15359_2757# a_15712_3988# 7.49e-21
C176 a_15868_2881# a_14791_2515# 1.46e-19
C177 a_15237_2515# a_15046_2515# 4.61e-19
C178 vd a_16024_5320# 0.0626f
C179 vd sensor_0.b 0.0693f
C180 a_14791_2515# a_15048_3988# 1.82e-19
C181 vpwr a_15815_2515# 7.93e-19
C182 a_14791_2515# a_15881_2489# 0.0426f
C183 a_15359_2757# a_15141_2515# 0.21f
C184 out_sigma out 5.44f
C185 sigma-delta_0.x1.D a_14791_2515# 0.229f
C186 a_14625_2515# a_15359_2757# 0.0701f
C187 buffer_0.d buffer_0.c 0.0518f
C188 out_buff a_15380_3988# 5.35e-19
C189 a_15380_3988# a_15214_5320# 0.00473f
C190 a_15712_3988# a_14716_3988# 2.04e-19
C191 a_16190_3988# a_15881_2489# 4.27e-19
C192 out_sigma a_16854_3988# 7.61e-19
C193 clk out_sigma 0.382f
C194 vd out 0.145p
C195 a_16024_5320# a_15712_3988# 0.00827f
C196 vpwr a_15359_2757# 0.378f
C197 sensor_0.d sensor_0.b 0.0152f
C198 sigma-delta_0.x1.Q a_16445_2515# 0.226f
C199 out_sigma a_15048_3988# 0.0146f
C200 a_15237_2515# a_15359_2757# 3.16e-19
C201 a_14625_2515# a_14716_3988# 1.47e-19
C202 buffer_0.a ib 0.00973f
C203 a_15546_5320# a_15380_3988# 0.00434f
C204 a_14882_5320# a_14716_3988# 0.00434f
C205 out_sigma a_14550_5320# 6.23e-19
C206 out_sigma a_15881_2489# 0.00735f
C207 a_15815_2515# a_15706_2515# 0.00742f
C208 vd a_16854_3988# 0.0174f
C209 clk vd 0.00542f
C210 sigma-delta_0.x1.D out_sigma 0.294f
C211 vpwr a_14716_3988# 0.0038f
C212 vd a_15048_3988# 0.00206f
C213 a_15359_2757# a_15403_2515# 3.69e-19
C214 out a_15712_3988# 0.18f
C215 vd a_14550_5320# 0.067f
C216 vd a_15881_2489# 0.00172f
C217 buffer_0.b out 0.00225f
C218 a_17020_5320# out 0.00192f
C219 a_16356_5320# a_16688_5320# 0.307f
C220 sigma-delta_0.x1.D vd 0.908f
C221 a_15359_2757# a_15706_2515# 0.0512f
C222 a_14791_2515# a_16445_2515# 2.01e-19
C223 a_15359_2757# a_15380_3988# 7.2e-20
C224 a_15712_3988# a_16854_3988# 0.00957f
C225 vd vts 0.94f
C226 out a_14882_5320# 0.0019f
C227 a_15249_2881# a_15141_2515# 0.0572f
C228 a_17020_5320# a_16854_3988# 0.00434f
C229 clk buffer_0.b 4.18e-19
C230 a_15868_2881# a_15712_3988# 5.54e-20
C231 a_15249_2881# a_14625_2515# 9.73e-19
C232 clk a_15141_2515# 3.26e-19
C233 a_16060_2515# clk 6.32e-21
C234 out_buff a_15214_5320# 5.44e-19
C235 a_15048_3988# a_15712_3988# 4.38e-19
C236 a_14625_2515# clk 0.274f
C237 a_15712_3988# a_15881_2489# 0.00381f
C238 sigma-delta_0.x1.D a_15712_3988# 0.339f
C239 out_sigma a_16445_2515# 0.0691f
C240 a_14625_2515# a_15048_3988# 1.92e-19
C241 vpwr a_15249_2881# 0.156f
C242 out_buff a_15546_5320# 2.84e-19
C243 a_16060_2515# a_15881_2489# 0.0074f
C244 a_15048_3988# a_14882_5320# 0.00482f
C245 a_16060_2515# sigma-delta_0.x1.D 4.54e-20
C246 a_14625_2515# a_15881_2489# 0.0436f
C247 sigma-delta_0.x1.D a_15141_2515# 0.00353f
C248 a_15546_5320# a_15214_5320# 0.296f
C249 vpwr clk 0.493f
C250 sensor_0.d vts 0.248f
C251 a_14882_5320# a_14550_5320# 0.296f
C252 a_15237_2515# clk 5.33e-20
C253 a_14625_2515# sigma-delta_0.x1.D 0.195f
C254 sensor_0.c sensor_0.b 0.55f
C255 buffer_0.b vts 0.112f
C256 a_15868_2881# vpwr 9.63e-19
C257 a_14791_2515# sigma-delta_0.x1.Q 0.00137f
C258 vpwr a_15048_3988# 0.00379f
C259 vd a_16445_2515# 0.00317f
C260 vpwr a_15881_2489# 0.688f
C261 a_16522_3988# a_16854_3988# 0.303f
C262 out_buff buffer_0.d 35.6f
C263 sensor_0.a sensor_0.b 0.821f
C264 vts buffer_0.c 0.416f
C265 vpwr sigma-delta_0.x1.D 0.483f
C266 sigma-delta_0.x1.Q a_16190_3988# 1.87e-20
C267 a_15237_2515# sigma-delta_0.x1.D 8.22e-19
C268 clk a_15403_2515# 1.82e-20
C269 ib vd 0.0124f
C270 buffer_0.a out_sigma 0.0182f
C271 a_16522_3988# a_15881_2489# 1.28e-20
C272 clk a_15706_2515# 6.46e-20
C273 a_16445_2515# a_15712_3988# 0.00366f
C274 a_15868_2881# a_15706_2515# 0.00645f
C275 sigma-delta_0.x1.Q out_sigma 0.668f
C276 sigma-delta_0.x1.D a_15403_2515# 5.41e-20
C277 out_buff a_14716_3988# 0.307f
C278 a_15048_3988# a_15380_3988# 0.302f
C279 buffer_0.a vd 5.58f
C280 a_16356_5320# a_16024_5320# 0.3f
C281 a_15706_2515# a_15881_2489# 0.251f
C282 a_15359_2757# a_15815_2515# 4.2e-19
C283 sigma-delta_0.x1.D a_15706_2515# 9.45e-19
C284 a_14625_2515# a_16445_2515# 4.71e-20
C285 out_buff a_16024_5320# 3.49e-20
C286 clk gnd 3.47f
C287 ib gnd 6.34f
C288 out_buff gnd 14.5f
C289 out gnd 59.9f
C290 out_sigma gnd 19.2f
C291 vpwr gnd 7.36f
C292 vts gnd 19.7f
C293 vd gnd 0.103p
C294 a_16060_2515# gnd 0.00223f
C295 a_15815_2515# gnd 9.68e-19
C296 a_15403_2515# gnd 0.00579f
C297 a_15237_2515# gnd 0.00863f
C298 a_15249_2881# gnd 0.00469f
C299 a_15046_2515# gnd 0.08f
C300 a_16445_2515# gnd 0.213f
C301 a_15706_2515# gnd 0.275f
C302 a_15881_2489# gnd 0.74f
C303 a_15141_2515# gnd 0.281f
C304 a_15359_2757# gnd 0.194f
C305 a_14791_2515# gnd 0.332f
C306 sigma-delta_0.x1.D gnd 2.56f
C307 a_14625_2515# gnd 0.7f
C308 sigma-delta_0.x1.Q gnd 1.09f
C309 a_17020_5320# gnd 0.557f
C310 a_16854_3988# gnd 0.348f
C311 a_16688_5320# gnd 0.388f
C312 a_16522_3988# gnd 0.356f
C313 a_16356_5320# gnd 0.392f
C314 a_16190_3988# gnd 0.357f
C315 a_16024_5320# gnd 0.447f
C316 a_15712_3988# gnd 69.7f
C317 a_15546_5320# gnd 0.449f
C318 a_15380_3988# gnd 0.365f
C319 a_15214_5320# gnd 0.387f
C320 a_15048_3988# gnd 0.364f
C321 a_14882_5320# gnd 0.39f
C322 a_14716_3988# gnd 0.366f
C323 a_14550_5320# gnd 0.587f
C324 buffer_0.c gnd 1.15f
C325 buffer_0.b gnd 2.31f
C326 buffer_0.a gnd 2.47f
C327 buffer_0.d gnd 20.1f
C328 sensor_0.b gnd 16.7f
C329 sensor_0.c gnd 0.658f
C330 sensor_0.a gnd 5.59f
C331 sensor_0.d gnd 0.293f
C332 a_6126_29386# gnd 0.593f
C333 out.t0 gnd 0.0079f
C334 out.t3 gnd 13.1f
C335 out.t2 gnd 28.9f
C336 out.t1 gnd 19.8f
C337 out.n0 gnd 10.6f
C338 out.n1 gnd 16.3f
C339 out.n2 gnd 61.4f
C340 out_sigma.t1 gnd 0.0149f
C341 out_sigma.t0 gnd 0.011f
C342 out_sigma.n0 gnd 0.245f
C343 out_sigma.t2 gnd 0.0325f
C344 out_sigma.n1 gnd 2.85f
C345 out_sigma.n2 gnd 1.76f
C346 vts.t17 gnd 0.1f
C347 vts.t20 gnd 0.00611f
C348 vts.t6 gnd 0.00573f
C349 vts.t3 gnd 0.00573f
C350 vts.n0 gnd 0.0271f
C351 vts.t1 gnd 0.00573f
C352 vts.t16 gnd 0.00573f
C353 vts.n1 gnd 0.0271f
C354 vts.t14 gnd 0.00573f
C355 vts.t12 gnd 0.00573f
C356 vts.n2 gnd 0.0271f
C357 vts.t10 gnd 0.00573f
C358 vts.t8 gnd 0.00573f
C359 vts.n3 gnd 0.0271f
C360 vts.t23 gnd 0.00616f
C361 vts.t21 gnd 0.1f
C362 vts.t24 gnd 0.00603f
C363 vts.n4 gnd 0.12f
C364 vts.n5 gnd 0.0685f
C365 vts.n6 gnd 0.0461f
C366 vts.n7 gnd 0.0538f
C367 vts.n8 gnd 0.0538f
C368 vts.n9 gnd 0.0457f
C369 vts.n10 gnd 0.0683f
C370 vts.n11 gnd 0.0645f
C371 vts.t19 gnd 0.0061f
C372 vts.n12 gnd 0.0548f
C373 vts.n13 gnd 0.00516f
C374 vts.n14 gnd 0.00536f
C375 vts.n15 gnd 0.0344f
C376 vts.n16 gnd 0.0344f
C377 vts.t2 gnd 0.272f
C378 vts.t5 gnd 0.333f
C379 vts.t18 gnd 0.337f
C380 vts.t22 gnd 0.355f
C381 vts.n17 gnd 0.279f
C382 vts.n18 gnd 0.0688f
C383 vts.t0 gnd 0.272f
C384 vts.t15 gnd 0.213f
C385 vts.t7 gnd 0.336f
C386 vts.t9 gnd 0.272f
C387 vts.t11 gnd 0.272f
C388 vts.t13 gnd 0.195f
C389 vts.n19 gnd 0.0653f
C390 vts.n20 gnd 0.0653f
C391 vts.n21 gnd 0.136f
C392 vts.n22 gnd 0.0628f
C393 vts.n23 gnd 0.0628f
C394 vts.n24 gnd 0.0317f
C395 vts.n25 gnd 0.032f
C396 vts.n26 gnd 0.196f
C397 vts.n28 gnd 0.00534f
C398 vts.n29 gnd 0.0103f
C399 vts.n30 gnd 0.00449f
C400 vts.t4 gnd 0.0378f
C401 vts.n31 gnd 0.342f
C402 vts.n32 gnd 8.23e-19
C403 vts.n33 gnd 0.002f
C404 vts.n34 gnd 0.0346f
C405 vts.t25 gnd 0.0138f
C406 vts.n35 gnd 0.669f
C407 vts.n36 gnd 0.833f
C408 buffer_0.d.n0 gnd 0.621f
C409 buffer_0.d.n1 gnd 0.584f
C410 buffer_0.d.t12 gnd 0.274f
C411 buffer_0.d.t13 gnd 0.274f
C412 buffer_0.d.n2 gnd 0.241f
C413 buffer_0.d.t9 gnd 0.274f
C414 buffer_0.d.n3 gnd 0.121f
C415 buffer_0.d.t7 gnd 0.274f
C416 buffer_0.d.n4 gnd 0.149f
C417 buffer_0.d.t11 gnd 33f
C418 buffer_0.d.n5 gnd 0.272f
C419 buffer_0.d.t10 gnd 0.021f
C420 buffer_0.d.t8 gnd 0.021f
C421 buffer_0.d.n6 gnd 0.112f
C422 buffer_0.d.n7 gnd 0.229f
C423 buffer_0.d.t2 gnd 0.701f
C424 buffer_0.d.n8 gnd 0.309f
C425 buffer_0.d.t1 gnd 0.0632f
C426 buffer_0.d.t3 gnd 0.434f
C427 buffer_0.d.t4 gnd 0.701f
C428 buffer_0.d.n9 gnd 0.309f
C429 buffer_0.d.t0 gnd 0.0631f
C430 buffer_0.d.t5 gnd 0.0631f
C431 buffer_0.d.t6 gnd 0.367f
C432 vtd.n0 gnd 0.544f
C433 vtd.n1 gnd 0.544f
C434 vtd.n2 gnd 0.544f
C435 vtd.n3 gnd 0.957f
C436 vtd.n4 gnd 0.174f
C437 vtd.n5 gnd 0.234f
C438 vtd.n6 gnd 0.321f
C439 vtd.t25 gnd 2.06f
C440 vtd.t29 gnd 0.402f
C441 vtd.n7 gnd 1.26f
C442 vtd.t27 gnd 0.401f
C443 vtd.t28 gnd 0.398f
C444 vtd.n8 gnd 0.396f
C445 vtd.t26 gnd 0.398f
C446 vtd.n9 gnd 0.204f
C447 vtd.t24 gnd 0.398f
C448 vtd.t1 gnd 0.0204f
C449 vtd.t5 gnd 0.0115f
C450 vtd.n10 gnd 0.436f
C451 vtd.t2 gnd 0.0115f
C452 vtd.n11 gnd 0.235f
C453 vtd.t6 gnd 0.0114f
C454 vtd.n12 gnd 0.247f
C455 vtd.t3 gnd 0.0114f
C456 vtd.t0 gnd 0.0115f
C457 vtd.t4 gnd 0.0205f
C458 vtd.n13 gnd 0.398f
C459 vtd.t7 gnd 0.0114f
C460 vtd.n14 gnd 0.218f
C461 vtd.n15 gnd 0.322f
C462 vtd.n16 gnd 0.45f
C463 vtd.t11 gnd 0.0239f
C464 vtd.t10 gnd 0.398f
C465 vtd.t20 gnd 0.398f
C466 vtd.t21 gnd 0.0228f
C467 vtd.t19 gnd 0.0228f
C468 vtd.t18 gnd 0.398f
C469 vtd.t12 gnd 0.398f
C470 vtd.t13 gnd 0.0228f
C471 vtd.t9 gnd 0.0228f
C472 vtd.t8 gnd 0.398f
C473 vtd.t22 gnd 0.398f
C474 vtd.t23 gnd 0.0228f
C475 vtd.t17 gnd 0.0228f
C476 vtd.t16 gnd 0.398f
C477 vtd.t14 gnd 0.398f
C478 vtd.t15 gnd 0.0237f
C479 vtd.n17 gnd 0.529f
C480 vtd.n18 gnd 0.339f
C481 vtd.n19 gnd 0.339f
C482 vtd.n20 gnd 0.622f
C483 vpwr.n0 gnd 7.54e-19
C484 vpwr.n1 gnd 5.58e-19
C485 vpwr.n2 gnd 0.00129f
C486 vpwr.t22 gnd 0.00331f
C487 vpwr.n3 gnd 0.00192f
C488 vpwr.n4 gnd 0.00211f
C489 vpwr.n5 gnd 8.86e-19
C490 vpwr.t31 gnd 0.00204f
C491 vpwr.n6 gnd 0.00253f
C492 vpwr.n7 gnd 0.00412f
C493 vpwr.n8 gnd 5.25e-19
C494 vpwr.n9 gnd 5.58e-19
C495 vpwr.n10 gnd 5.58e-19
C496 vpwr.n11 gnd 0.00129f
C497 vpwr.n12 gnd 0.00855f
C498 vpwr.n13 gnd 5.92e-19
C499 vpwr.t30 gnd 0.00155f
C500 vpwr.t25 gnd 0.00391f
C501 vpwr.n14 gnd 0.00669f
C502 vpwr.n15 gnd 0.00264f
C503 vpwr.n16 gnd 0.00193f
C504 vpwr.n17 gnd 3.77e-19
C505 vpwr.n18 gnd 3.47e-19
C506 vpwr.n19 gnd 7.75e-19
C507 vpwr.n20 gnd 0.00273f
C508 vpwr.n21 gnd 5.32e-19
C509 vpwr.n22 gnd 0.00261f
C510 vpwr.n23 gnd 6.22e-19
C511 vpwr.n24 gnd 7.41e-19
C512 vpwr.n25 gnd 0.00193f
C513 vpwr.n26 gnd 0.0404f
C514 vpwr.n27 gnd 0.0636f
C515 vpwr.n28 gnd 0.492f
C516 vpwr.n29 gnd 0.0803f
C517 vpwr.n30 gnd 0.00889f
C518 vpwr.t18 gnd 0.00153f
C519 vpwr.t13 gnd 0.00153f
C520 vpwr.n31 gnd 0.00331f
C521 vpwr.t21 gnd 0.00355f
C522 vpwr.n32 gnd 0.00793f
C523 vpwr.n33 gnd 0.00784f
C524 vpwr.n34 gnd 0.00163f
C525 vpwr.n35 gnd 0.00784f
C526 vpwr.n36 gnd 0.00784f
C527 vpwr.t7 gnd 0.00681f
C528 vpwr.n37 gnd 0.00278f
C529 vpwr.n38 gnd 0.00784f
C530 vpwr.t24 gnd 0.00101f
C531 vpwr.t3 gnd 0.0019f
C532 vpwr.n39 gnd 0.0031f
C533 vpwr.n40 gnd 0.0047f
C534 vpwr.t1 gnd 0.00228f
C535 vpwr.t11 gnd 0.00103f
C536 vpwr.n41 gnd 0.00896f
C537 vpwr.n42 gnd 0.0537f
C538 vpwr.t5 gnd 0.003f
C539 vpwr.t15 gnd 0.00108f
C540 vpwr.n43 gnd 0.00399f
C541 vpwr.n44 gnd 0.00707f
C542 vpwr.n45 gnd 0.00563f
C543 vpwr.n46 gnd 0.00381f
C544 vpwr.n47 gnd 0.0115f
C545 vpwr.n48 gnd 0.00784f
C546 vpwr.n49 gnd 0.00216f
C547 vpwr.n50 gnd 0.00741f
C548 vpwr.n51 gnd 0.0022f
C549 vpwr.n52 gnd 0.00784f
C550 vpwr.n53 gnd 0.00784f
C551 vpwr.n54 gnd 0.00784f
C552 vpwr.n55 gnd 0.00267f
C553 vpwr.n56 gnd 0.0109f
C554 vpwr.n57 gnd 0.00176f
C555 vpwr.t27 gnd 0.00101f
C556 vpwr.t29 gnd 0.00149f
C557 vpwr.n58 gnd 0.00269f
C558 vpwr.n59 gnd 0.00723f
C559 vpwr.n60 gnd 0.00154f
C560 vpwr.n61 gnd 0.00784f
C561 vpwr.n62 gnd 0.00784f
C562 vpwr.n63 gnd 0.00784f
C563 vpwr.n64 gnd 0.00278f
C564 vpwr.n65 gnd 0.00278f
C565 vpwr.n66 gnd 0.00268f
C566 vpwr.n67 gnd 0.00784f
C567 vpwr.n68 gnd 0.00784f
C568 vpwr.n69 gnd 0.00784f
C569 vpwr.n70 gnd 0.00211f
C570 vpwr.n71 gnd 0.00231f
C571 vpwr.n72 gnd 0.00978f
C572 vpwr.n73 gnd 0.00708f
C573 vpwr.n74 gnd 0.00695f
C574 vpwr.n75 gnd 0.00675f
C575 vpwr.t10 gnd 0.0545f
C576 vpwr.t0 gnd 0.045f
C577 vpwr.t4 gnd 0.0545f
C578 vpwr.t14 gnd 0.0353f
C579 vpwr.t23 gnd 0.0273f
C580 vpwr.t2 gnd 0.0273f
C581 vpwr.t9 gnd 0.0242f
C582 vpwr.t19 gnd 0.0263f
C583 vpwr.t6 gnd 0.0422f
C584 vpwr.t26 gnd 0.0419f
C585 vpwr.t28 gnd 0.0337f
C586 vpwr.t16 gnd 0.034f
C587 vpwr.t8 gnd 0.0272f
C588 vpwr.t20 gnd 0.0511f
C589 vpwr.t17 gnd 0.05f
C590 vpwr.t12 gnd 0.0219f
C591 vpwr.n76 gnd 0.00239f
C592 vpwr.n77 gnd 0.0593f
C593 vpwr.n78 gnd 0.00316f
C594 vpwr.n79 gnd 0.0012f
C595 vpwr.n80 gnd 0.00543f
C596 vpwr.n81 gnd 0.00177f
C597 vpwr.n82 gnd 0.00561f
C598 vpwr.n83 gnd 0.0366f
C599 vd.t74 gnd 21f
C600 vd.t75 gnd 21f
C601 vd.t73 gnd 41.7f
C602 vd.n0 gnd 20.8f
C603 vd.n1 gnd 13.3f
C604 vd.t46 gnd 0.0555f
C605 vd.n2 gnd 17f
C606 vd.n3 gnd 0.0138f
C607 vd.n4 gnd 0.00341f
C608 vd.n5 gnd 0.0104f
C609 vd.n6 gnd 6.53e-19
C610 vd.t1 gnd 0.00768f
C611 vd.n7 gnd 0.00182f
C612 vd.n8 gnd 0.012f
C613 vd.n9 gnd 0.00247f
C614 vd.n10 gnd 0.0138f
C615 vd.n11 gnd 7.06e-19
C616 vd.n12 gnd 0.00505f
C617 vd.n13 gnd 0.0138f
C618 vd.t0 gnd 0.145f
C619 vd.n15 gnd 0.0137f
C620 vd.n16 gnd 0.00505f
C621 vd.n18 gnd 0.139f
C622 vd.n19 gnd 0.0185f
C623 vd.n20 gnd 0.0137f
C624 vd.n21 gnd 0.00562f
C625 vd.n22 gnd 0.00929f
C626 vd.n23 gnd 0.121f
C627 vd.n24 gnd 0.00939f
C628 vd.n25 gnd 0.00574f
C629 vd.n26 gnd 0.0146f
C630 vd.n27 gnd 0.0293f
C631 vd.n28 gnd 0.0148f
C632 vd.n29 gnd 0.00811f
C633 vd.n30 gnd 0.0447f
C634 vd.n31 gnd 0.00317f
C635 vd.n32 gnd 0.00855f
C636 vd.n33 gnd 0.00176f
C637 vd.n34 gnd 0.00229f
C638 vd.n35 gnd 0.00212f
C639 vd.n36 gnd 0.0103f
C640 vd.n37 gnd 0.0136f
C641 vd.n38 gnd 0.131f
C642 vd.n39 gnd 0.0719f
C643 vd.n40 gnd 0.0539f
C644 vd.n41 gnd 0.0798f
C645 vd.n42 gnd 0.586f
C646 vd.t29 gnd -0.0168f
C647 vd.t47 gnd 0.786f
C648 vd.n43 gnd 0.098f
C649 vd.t10 gnd 0.582f
C650 vd.t40 gnd 0.758f
C651 vd.t8 gnd 0.61f
C652 vd.n44 gnd 0.397f
C653 vd.n45 gnd 0.0647f
C654 vd.n46 gnd 0.0647f
C655 vd.n47 gnd 0.0647f
C656 vd.t43 gnd 0.759f
C657 vd.t2 gnd 0.168f
C658 vd.t4 gnd 0.168f
C659 vd.t6 gnd 0.168f
C660 vd.t15 gnd 0.168f
C661 vd.t12 gnd 0.168f
C662 vd.t14 gnd 0.142f
C663 vd.n48 gnd 0.0679f
C664 vd.n49 gnd 0.0633f
C665 vd.t61 gnd 0.138f
C666 vd.t64 gnd 0.168f
C667 vd.t57 gnd 0.168f
C668 vd.t66 gnd 0.168f
C669 vd.t68 gnd 0.168f
C670 vd.t62 gnd 0.168f
C671 vd.t26 gnd -0.0179f
C672 vd.n50 gnd 0.0799f
C673 vd.t70 gnd 0.596f
C674 vd.n51 gnd 0.398f
C675 vd.t59 gnd 0.599f
C676 vd.t42 gnd 0.756f
C677 vd.n52 gnd 0.623f
C678 vd.n53 gnd 0.0979f
C679 vd.n54 gnd 0.169f
C680 vd.n55 gnd 0.505f
C681 vd.n56 gnd 0.0783f
C682 vd.n57 gnd 0.0783f
C683 vd.n58 gnd 0.098f
C684 vd.n59 gnd 0.0647f
C685 vd.n60 gnd 0.0793f
C686 vd.n61 gnd 0.0793f
C687 vd.n62 gnd 0.493f
C688 vd.n63 gnd 0.186f
C689 vd.n64 gnd 0.0985f
C690 vd.n65 gnd 0.0716f
C691 vd.n66 gnd 0.0654f
C692 vd.n67 gnd 0.00382f
C693 vd.t13 gnd 0.00256f
C694 vd.t16 gnd 0.00256f
C695 vd.n68 gnd 0.00876f
C696 vd.n69 gnd 0.0086f
C697 vd.t3 gnd 0.00256f
C698 vd.t30 gnd 0.00256f
C699 vd.n70 gnd 0.0116f
C700 vd.t28 gnd 0.0552f
C701 vd.t31 gnd 0.00263f
C702 vd.n71 gnd 0.0814f
C703 vd.n72 gnd 0.022f
C704 vd.t7 gnd 0.00256f
C705 vd.t5 gnd 0.00256f
C706 vd.n73 gnd 0.0143f
C707 vd.n74 gnd 0.0189f
C708 vd.n75 gnd 0.0104f
C709 vd.n76 gnd 0.00127f
C710 vd.n77 gnd 0.0116f
C711 vd.t11 gnd 0.0384f
C712 vd.t9 gnd 0.0384f
C713 vd.n78 gnd 0.324f
C714 vd.n79 gnd 0.271f
C715 vd.t60 gnd 0.0384f
C716 vd.t71 gnd 0.0384f
C717 vd.n80 gnd 0.347f
C718 vd.t25 gnd 0.0552f
C719 vd.n81 gnd 0.0882f
C720 vd.t27 gnd 0.00525f
C721 vd.t63 gnd 0.00256f
C722 vd.n82 gnd 0.0123f
C723 vd.n83 gnd 0.0129f
C724 vd.t69 gnd 0.00256f
C725 vd.t67 gnd 0.00256f
C726 vd.n84 gnd 0.0143f
C727 vd.n85 gnd 0.0196f
C728 vd.t58 gnd 0.00256f
C729 vd.t65 gnd 0.00256f
C730 vd.n86 gnd 0.0105f
C731 vd.n87 gnd 0.0389f
C732 vd.n88 gnd 0.23f
C733 vd.n89 gnd 0.057f
C734 vd.n90 gnd 0.00405f
C735 vd.n91 gnd 1.23f
C736 vd.t34 gnd 0.00512f
C737 vd.t32 gnd 0.0896f
C738 vd.t35 gnd 0.00512f
C739 vd.t37 gnd 0.00574f
C740 vd.n92 gnd 0.0865f
C741 vd.n93 gnd 0.072f
C742 vd.n94 gnd 0.0922f
C743 vd.n95 gnd 0.0558f
C744 vd.n96 gnd 0.282f
C745 vd.n97 gnd 0.225f
C746 vd.n98 gnd 0.0184f
C747 vd.n99 gnd 0.0184f
C748 vd.t41 gnd 0.0911f
C749 vd.t33 gnd 0.0984f
C750 vd.t38 gnd 0.338f
C751 vd.n100 gnd 0.269f
C752 vd.n101 gnd 0.0105f
C753 vd.t48 gnd 0.151f
C754 vd.n102 gnd 0.19f
C755 vd.n103 gnd 0.0138f
C756 vd.n104 gnd 0.0136f
C757 vd.n105 gnd 0.0115f
C758 vd.t21 gnd 0.0897f
C759 vd.t45 gnd 0.00594f
C760 vd.t23 gnd 0.00512f
C761 vd.n106 gnd 0.0839f
C762 vd.n107 gnd 0.0687f
C763 vd.t24 gnd 0.00512f
C764 vd.n108 gnd 0.0728f
C765 vd.n109 gnd 0.00171f
C766 vd.t20 gnd 0.00512f
C767 vd.n110 gnd 0.0297f
C768 vd.t19 gnd 0.00539f
C769 vd.t54 gnd 0.00511f
C770 vd.t56 gnd 0.00511f
C771 vd.n111 gnd 0.0406f
C772 vd.n112 gnd 0.0527f
C773 vd.t17 gnd 0.0895f
C774 vd.n113 gnd 0.0593f
C775 vd.n114 gnd 0.00602f
C776 vd.n115 gnd 0.00276f
C777 vd.n116 gnd 0.0493f
C778 vd.n117 gnd 0.0574f
C779 vd.n118 gnd 0.337f
C780 vd.t18 gnd 0.228f
C781 vd.n119 gnd 0.279f
C782 vd.n120 gnd 0.0217f
C783 vd.n121 gnd 0.0216f
C784 vd.t53 gnd 0.411f
C785 vd.t55 gnd 0.256f
C786 vd.n122 gnd 0.19f
C787 vd.n123 gnd 0.0136f
C788 vd.n124 gnd 0.0147f
C789 vd.n125 gnd 0.115f
C790 vd.n126 gnd 0.139f
C791 vd.t49 gnd 0.0999f
C792 vd.t44 gnd 0.0793f
C793 vd.n127 gnd 0.0819f
C794 vd.n128 gnd 0.0819f
C795 vd.n129 gnd 0.165f
C796 vd.n130 gnd 0.00585f
C797 vd.n131 gnd 0.00583f
C798 vd.t51 gnd 0.244f
C799 vd.n132 gnd 0.281f
C800 vd.n133 gnd 0.0168f
C801 vd.n134 gnd 0.0165f
C802 vd.t50 gnd 0.132f
C803 vd.t52 gnd 0.264f
C804 vd.t22 gnd 0.167f
C805 vd.n135 gnd 0.115f
C806 vd.n136 gnd 0.0111f
C807 vd.n137 gnd 0.0121f
C808 vd.n138 gnd 0.113f
C809 vd.n139 gnd 0.284f
C810 vd.n140 gnd 0.009f
C811 vd.n141 gnd 0.00889f
C812 vd.t36 gnd 0.19f
C813 vd.t39 gnd 0.187f
C814 vd.t72 gnd 0.287f
C815 vd.n142 gnd 0.19f
C816 vd.n143 gnd 0.0127f
C817 vd.n144 gnd 0.0138f
C818 vd.n145 gnd 0.161f
C819 vd.n146 gnd 0.0931f
C820 vd.n147 gnd 0.547f
C821 vd.n148 gnd 5.86f
C822 vd.n149 gnd 4.83f
C823 vd.n150 gnd 0.446f
C824 out_buff.t6 gnd 0.0642f
C825 out_buff.t2 gnd 0.308f
C826 out_buff.t9 gnd 0.0461f
C827 out_buff.n0 gnd 0.17f
C828 out_buff.t1 gnd 0.511f
C829 out_buff.n1 gnd 0.235f
C830 out_buff.n2 gnd 0.051f
C831 out_buff.t5 gnd 0.264f
C832 out_buff.t8 gnd 0.0461f
C833 out_buff.t4 gnd 0.0461f
C834 out_buff.n3 gnd 0.17f
C835 out_buff.t3 gnd 0.511f
C836 out_buff.n4 gnd 0.234f
C837 out_buff.n5 gnd 0.0511f
C838 out_buff.t11 gnd 0.0103f
C839 out_buff.t10 gnd 38.6f
C840 out_buff.n6 gnd 0.465f
C841 out_buff.t0 gnd 0.0154f
C842 out_buff.t7 gnd 0.0154f
C843 out_buff.n7 gnd 0.111f
C844 out_buff.n8 gnd 0.0709f
C845 out_buff.n9 gnd 0.223f
C846 out_buff.n10 gnd 0.225f
C847 out_buff.n11 gnd 0.495f
C848 out_buff.n12 gnd 1.31f
C849 out_buff.n13 gnd 0.256f
C850 buffer_0.b.n0 gnd 0.0408f
C851 buffer_0.b.n1 gnd 0.0786f
C852 buffer_0.b.t8 gnd 0.0101f
C853 buffer_0.b.t6 gnd 0.0101f
C854 buffer_0.b.n2 gnd 0.0936f
C855 buffer_0.b.t4 gnd 0.0101f
C856 buffer_0.b.t2 gnd 0.0101f
C857 buffer_0.b.n3 gnd 0.0563f
C858 buffer_0.b.n4 gnd 0.0779f
C859 buffer_0.b.n5 gnd 0.0463f
C860 buffer_0.b.t17 gnd 1.68f
C861 buffer_0.b.t16 gnd 1.67f
C862 buffer_0.b.n6 gnd 1.6f
C863 buffer_0.b.t7 gnd 0.126f
C864 buffer_0.b.t5 gnd 0.202f
C865 buffer_0.b.n7 gnd 0.291f
C866 buffer_0.b.t3 gnd 0.202f
C867 buffer_0.b.n8 gnd 0.16f
C868 buffer_0.b.t1 gnd 0.202f
C869 buffer_0.b.n9 gnd 0.16f
C870 buffer_0.b.t14 gnd 0.202f
C871 buffer_0.b.n10 gnd 0.163f
C872 buffer_0.b.t11 gnd 0.202f
C873 buffer_0.b.t13 gnd 0.0104f
C874 buffer_0.b.n11 gnd 0.324f
C875 buffer_0.b.n12 gnd 0.00756f
C876 buffer_0.b.n13 gnd 0.00153f
C877 buffer_0.b.t15 gnd 0.0101f
C878 buffer_0.b.t12 gnd 0.0101f
C879 buffer_0.b.n14 gnd 0.0684f
C880 buffer_0.b.t9 gnd 0.024f
C881 buffer_0.b.t0 gnd 0.0172f
C882 buffer_0.b.t10 gnd 0.0356f
C883 buffer_0.b.n15 gnd 0.224f
C884 buffer_0.b.n16 gnd 0.161f
C885 sensor_0.a.n0 gnd 0.396f
C886 sensor_0.a.n1 gnd 0.413f
C887 sensor_0.a.t15 gnd 0.277f
C888 sensor_0.a.t14 gnd 0.276f
C889 sensor_0.a.n2 gnd 0.293f
C890 sensor_0.a.t12 gnd 0.276f
C891 sensor_0.a.n3 gnd 0.15f
C892 sensor_0.a.t13 gnd 0.276f
C893 sensor_0.a.n4 gnd 0.148f
C894 sensor_0.a.t9 gnd 0.0159f
C895 sensor_0.a.t8 gnd 0.276f
C896 sensor_0.a.t10 gnd 0.276f
C897 sensor_0.a.t11 gnd 0.0177f
C898 sensor_0.a.t7 gnd 0.0141f
C899 sensor_0.a.t4 gnd 0.00791f
C900 sensor_0.a.n5 gnd 0.277f
C901 sensor_0.a.t3 gnd 0.00792f
C902 sensor_0.a.n6 gnd 0.152f
C903 sensor_0.a.t0 gnd 0.00792f
C904 sensor_0.a.n7 gnd 0.19f
C905 sensor_0.a.t2 gnd 0.0141f
C906 sensor_0.a.t6 gnd 0.00791f
C907 sensor_0.a.n8 gnd 0.276f
C908 sensor_0.a.t1 gnd 0.0079f
C909 sensor_0.a.n9 gnd 0.154f
C910 sensor_0.a.t5 gnd 0.00792f
C911 sensor_0.a.n10 gnd 0.19f
C912 sensor_0.a.n11 gnd 0.384f
C913 sensor_0.b.t16 gnd 0.0077f
C914 sensor_0.b.t18 gnd 0.0077f
C915 sensor_0.b.n0 gnd 0.0683f
C916 sensor_0.b.t17 gnd 0.0077f
C917 sensor_0.b.t19 gnd 0.0077f
C918 sensor_0.b.n1 gnd 0.0506f
C919 sensor_0.b.n2 gnd 0.162f
C920 sensor_0.b.t3 gnd 0.00651f
C921 sensor_0.b.t11 gnd 0.00386f
C922 sensor_0.b.n3 gnd 0.139f
C923 sensor_0.b.t5 gnd 0.00385f
C924 sensor_0.b.n4 gnd 0.0928f
C925 sensor_0.b.t13 gnd 0.00385f
C926 sensor_0.b.n5 gnd 0.137f
C927 sensor_0.b.n6 gnd 0.202f
C928 sensor_0.b.t2 gnd 0.134f
C929 sensor_0.b.t10 gnd 0.127f
C930 sensor_0.b.t4 gnd 0.127f
C931 sensor_0.b.t12 gnd 0.0845f
C932 sensor_0.b.t32 gnd 0.134f
C933 sensor_0.b.t24 gnd 0.127f
C934 sensor_0.b.t31 gnd 0.127f
C935 sensor_0.b.t23 gnd 0.0845f
C936 sensor_0.b.t26 gnd 0.134f
C937 sensor_0.b.t34 gnd 0.127f
C938 sensor_0.b.t21 gnd 0.127f
C939 sensor_0.b.t29 gnd 0.0845f
C940 sensor_0.b.t20 gnd 0.134f
C941 sensor_0.b.t27 gnd 0.127f
C942 sensor_0.b.t28 gnd 0.127f
C943 sensor_0.b.t35 gnd 0.0845f
C944 sensor_0.b.t30 gnd 0.134f
C945 sensor_0.b.t22 gnd 0.127f
C946 sensor_0.b.t33 gnd 0.127f
C947 sensor_0.b.t25 gnd 0.0856f
C948 sensor_0.b.n7 gnd 0.119f
C949 sensor_0.b.n8 gnd 0.0626f
C950 sensor_0.b.n9 gnd 0.0626f
C951 sensor_0.b.n10 gnd 0.0626f
C952 sensor_0.b.t0 gnd 0.134f
C953 sensor_0.b.t8 gnd 0.127f
C954 sensor_0.b.t6 gnd 0.127f
C955 sensor_0.b.t14 gnd 0.0845f
C956 sensor_0.b.n11 gnd 0.0519f
C957 sensor_0.b.t1 gnd 0.00705f
C958 sensor_0.b.t9 gnd 0.00386f
C959 sensor_0.b.n12 gnd 0.138f
C960 sensor_0.b.t7 gnd 0.00386f
C961 sensor_0.b.n13 gnd 0.073f
C962 sensor_0.b.t15 gnd 0.00389f
C963 sensor_0.b.n14 gnd 0.0704f
C964 sensor_0.b.n15 gnd 0.0509f
C965 buffer_0.a.n0 gnd 0.146f
C966 buffer_0.a.t2 gnd 0.149f
C967 buffer_0.a.n1 gnd 0.323f
C968 buffer_0.a.t3 gnd 0.014f
C969 buffer_0.a.t12 gnd 0.00689f
C970 buffer_0.a.n2 gnd 0.0272f
C971 buffer_0.a.t11 gnd 0.149f
C972 buffer_0.a.t14 gnd 0.00689f
C973 buffer_0.a.t1 gnd 0.00689f
C974 buffer_0.a.n3 gnd 0.0627f
C975 buffer_0.a.t10 gnd 0.00689f
C976 buffer_0.a.t8 gnd 0.00689f
C977 buffer_0.a.n4 gnd 0.0384f
C978 buffer_0.a.n5 gnd 0.0492f
C979 buffer_0.a.t9 gnd 0.149f
C980 buffer_0.a.t7 gnd 0.149f
C981 buffer_0.a.t13 gnd 0.149f
C982 buffer_0.a.t16 gnd 1.15f
C983 buffer_0.a.t17 gnd 1.15f
C984 buffer_0.a.n6 gnd 0.98f
C985 buffer_0.a.t0 gnd 0.0876f
C986 buffer_0.a.n7 gnd 0.191f
C987 buffer_0.a.n8 gnd 0.0985f
C988 buffer_0.a.n9 gnd 0.0982f
C989 buffer_0.a.n10 gnd 0.026f
C990 buffer_0.a.n11 gnd 0.112f
C991 buffer_0.a.n12 gnd 0.00975f
C992 buffer_0.a.t15 gnd 0.0118f
C993 buffer_0.a.t5 gnd 0.0118f
C994 buffer_0.a.t4 gnd 0.0164f
C995 buffer_0.a.t6 gnd 0.0118f
C996 buffer_0.a.n13 gnd 0.136f
*.ends



**** end user architecture code
x1 vd out l0
.ends


* expanding   symbol:  /foss/designs/temp-sensor/ask_modulator/xschem/l0.sym # of pins=2
** sym_path: /foss/designs/temp-sensor/ask_modulator/xschem/l0.sym
** sch_path: /foss/designs/temp-sensor/ask_modulator/xschem/l0.sch
.subckt l0 p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 993p m=1
Cs1 p1 net1 58.53f m=1
Cs2 p2 net2 52.93f m=1
Rs1 net1 GND 24.1 m=1
Rs2 net2 GND 22.94 m=1
R1 p2 net3 3.443 m=1
.ends

.GLOBAL GND
.end
