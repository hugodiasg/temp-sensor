magic
tech sky130A
magscale 1 2
timestamp 1675569099
<< metal4 >>
rect -2309 53839 2309 53880
rect -2309 49841 2053 53839
rect 2289 49841 2309 53839
rect -2309 49800 2309 49841
rect -2309 49519 2309 49560
rect -2309 45521 2053 49519
rect 2289 45521 2309 49519
rect -2309 45480 2309 45521
rect -2309 45199 2309 45240
rect -2309 41201 2053 45199
rect 2289 41201 2309 45199
rect -2309 41160 2309 41201
rect -2309 40879 2309 40920
rect -2309 36881 2053 40879
rect 2289 36881 2309 40879
rect -2309 36840 2309 36881
rect -2309 36559 2309 36600
rect -2309 32561 2053 36559
rect 2289 32561 2309 36559
rect -2309 32520 2309 32561
rect -2309 32239 2309 32280
rect -2309 28241 2053 32239
rect 2289 28241 2309 32239
rect -2309 28200 2309 28241
rect -2309 27919 2309 27960
rect -2309 23921 2053 27919
rect 2289 23921 2309 27919
rect -2309 23880 2309 23921
rect -2309 23599 2309 23640
rect -2309 19601 2053 23599
rect 2289 19601 2309 23599
rect -2309 19560 2309 19601
rect -2309 19279 2309 19320
rect -2309 15281 2053 19279
rect 2289 15281 2309 19279
rect -2309 15240 2309 15281
rect -2309 14959 2309 15000
rect -2309 10961 2053 14959
rect 2289 10961 2309 14959
rect -2309 10920 2309 10961
rect -2309 10639 2309 10680
rect -2309 6641 2053 10639
rect 2289 6641 2309 10639
rect -2309 6600 2309 6641
rect -2309 6319 2309 6360
rect -2309 2321 2053 6319
rect 2289 2321 2309 6319
rect -2309 2280 2309 2321
rect -2309 1999 2309 2040
rect -2309 -1999 2053 1999
rect 2289 -1999 2309 1999
rect -2309 -2040 2309 -1999
rect -2309 -2321 2309 -2280
rect -2309 -6319 2053 -2321
rect 2289 -6319 2309 -2321
rect -2309 -6360 2309 -6319
rect -2309 -6641 2309 -6600
rect -2309 -10639 2053 -6641
rect 2289 -10639 2309 -6641
rect -2309 -10680 2309 -10639
rect -2309 -10961 2309 -10920
rect -2309 -14959 2053 -10961
rect 2289 -14959 2309 -10961
rect -2309 -15000 2309 -14959
rect -2309 -15281 2309 -15240
rect -2309 -19279 2053 -15281
rect 2289 -19279 2309 -15281
rect -2309 -19320 2309 -19279
rect -2309 -19601 2309 -19560
rect -2309 -23599 2053 -19601
rect 2289 -23599 2309 -19601
rect -2309 -23640 2309 -23599
rect -2309 -23921 2309 -23880
rect -2309 -27919 2053 -23921
rect 2289 -27919 2309 -23921
rect -2309 -27960 2309 -27919
rect -2309 -28241 2309 -28200
rect -2309 -32239 2053 -28241
rect 2289 -32239 2309 -28241
rect -2309 -32280 2309 -32239
rect -2309 -32561 2309 -32520
rect -2309 -36559 2053 -32561
rect 2289 -36559 2309 -32561
rect -2309 -36600 2309 -36559
rect -2309 -36881 2309 -36840
rect -2309 -40879 2053 -36881
rect 2289 -40879 2309 -36881
rect -2309 -40920 2309 -40879
rect -2309 -41201 2309 -41160
rect -2309 -45199 2053 -41201
rect 2289 -45199 2309 -41201
rect -2309 -45240 2309 -45199
rect -2309 -45521 2309 -45480
rect -2309 -49519 2053 -45521
rect 2289 -49519 2309 -45521
rect -2309 -49560 2309 -49519
rect -2309 -49841 2309 -49800
rect -2309 -53839 2053 -49841
rect 2289 -53839 2309 -49841
rect -2309 -53880 2309 -53839
<< via4 >>
rect 2053 49841 2289 53839
rect 2053 45521 2289 49519
rect 2053 41201 2289 45199
rect 2053 36881 2289 40879
rect 2053 32561 2289 36559
rect 2053 28241 2289 32239
rect 2053 23921 2289 27919
rect 2053 19601 2289 23599
rect 2053 15281 2289 19279
rect 2053 10961 2289 14959
rect 2053 6641 2289 10639
rect 2053 2321 2289 6319
rect 2053 -1999 2289 1999
rect 2053 -6319 2289 -2321
rect 2053 -10639 2289 -6641
rect 2053 -14959 2289 -10961
rect 2053 -19279 2289 -15281
rect 2053 -23599 2289 -19601
rect 2053 -27919 2289 -23921
rect 2053 -32239 2289 -28241
rect 2053 -36559 2289 -32561
rect 2053 -40879 2289 -36881
rect 2053 -45199 2289 -41201
rect 2053 -49519 2289 -45521
rect 2053 -53839 2289 -49841
<< mimcap2 >>
rect -2229 53760 1691 53800
rect -2229 49920 -2189 53760
rect 1651 49920 1691 53760
rect -2229 49880 1691 49920
rect -2229 49440 1691 49480
rect -2229 45600 -2189 49440
rect 1651 45600 1691 49440
rect -2229 45560 1691 45600
rect -2229 45120 1691 45160
rect -2229 41280 -2189 45120
rect 1651 41280 1691 45120
rect -2229 41240 1691 41280
rect -2229 40800 1691 40840
rect -2229 36960 -2189 40800
rect 1651 36960 1691 40800
rect -2229 36920 1691 36960
rect -2229 36480 1691 36520
rect -2229 32640 -2189 36480
rect 1651 32640 1691 36480
rect -2229 32600 1691 32640
rect -2229 32160 1691 32200
rect -2229 28320 -2189 32160
rect 1651 28320 1691 32160
rect -2229 28280 1691 28320
rect -2229 27840 1691 27880
rect -2229 24000 -2189 27840
rect 1651 24000 1691 27840
rect -2229 23960 1691 24000
rect -2229 23520 1691 23560
rect -2229 19680 -2189 23520
rect 1651 19680 1691 23520
rect -2229 19640 1691 19680
rect -2229 19200 1691 19240
rect -2229 15360 -2189 19200
rect 1651 15360 1691 19200
rect -2229 15320 1691 15360
rect -2229 14880 1691 14920
rect -2229 11040 -2189 14880
rect 1651 11040 1691 14880
rect -2229 11000 1691 11040
rect -2229 10560 1691 10600
rect -2229 6720 -2189 10560
rect 1651 6720 1691 10560
rect -2229 6680 1691 6720
rect -2229 6240 1691 6280
rect -2229 2400 -2189 6240
rect 1651 2400 1691 6240
rect -2229 2360 1691 2400
rect -2229 1920 1691 1960
rect -2229 -1920 -2189 1920
rect 1651 -1920 1691 1920
rect -2229 -1960 1691 -1920
rect -2229 -2400 1691 -2360
rect -2229 -6240 -2189 -2400
rect 1651 -6240 1691 -2400
rect -2229 -6280 1691 -6240
rect -2229 -6720 1691 -6680
rect -2229 -10560 -2189 -6720
rect 1651 -10560 1691 -6720
rect -2229 -10600 1691 -10560
rect -2229 -11040 1691 -11000
rect -2229 -14880 -2189 -11040
rect 1651 -14880 1691 -11040
rect -2229 -14920 1691 -14880
rect -2229 -15360 1691 -15320
rect -2229 -19200 -2189 -15360
rect 1651 -19200 1691 -15360
rect -2229 -19240 1691 -19200
rect -2229 -19680 1691 -19640
rect -2229 -23520 -2189 -19680
rect 1651 -23520 1691 -19680
rect -2229 -23560 1691 -23520
rect -2229 -24000 1691 -23960
rect -2229 -27840 -2189 -24000
rect 1651 -27840 1691 -24000
rect -2229 -27880 1691 -27840
rect -2229 -28320 1691 -28280
rect -2229 -32160 -2189 -28320
rect 1651 -32160 1691 -28320
rect -2229 -32200 1691 -32160
rect -2229 -32640 1691 -32600
rect -2229 -36480 -2189 -32640
rect 1651 -36480 1691 -32640
rect -2229 -36520 1691 -36480
rect -2229 -36960 1691 -36920
rect -2229 -40800 -2189 -36960
rect 1651 -40800 1691 -36960
rect -2229 -40840 1691 -40800
rect -2229 -41280 1691 -41240
rect -2229 -45120 -2189 -41280
rect 1651 -45120 1691 -41280
rect -2229 -45160 1691 -45120
rect -2229 -45600 1691 -45560
rect -2229 -49440 -2189 -45600
rect 1651 -49440 1691 -45600
rect -2229 -49480 1691 -49440
rect -2229 -49920 1691 -49880
rect -2229 -53760 -2189 -49920
rect 1651 -53760 1691 -49920
rect -2229 -53800 1691 -53760
<< mimcap2contact >>
rect -2189 49920 1651 53760
rect -2189 45600 1651 49440
rect -2189 41280 1651 45120
rect -2189 36960 1651 40800
rect -2189 32640 1651 36480
rect -2189 28320 1651 32160
rect -2189 24000 1651 27840
rect -2189 19680 1651 23520
rect -2189 15360 1651 19200
rect -2189 11040 1651 14880
rect -2189 6720 1651 10560
rect -2189 2400 1651 6240
rect -2189 -1920 1651 1920
rect -2189 -6240 1651 -2400
rect -2189 -10560 1651 -6720
rect -2189 -14880 1651 -11040
rect -2189 -19200 1651 -15360
rect -2189 -23520 1651 -19680
rect -2189 -27840 1651 -24000
rect -2189 -32160 1651 -28320
rect -2189 -36480 1651 -32640
rect -2189 -40800 1651 -36960
rect -2189 -45120 1651 -41280
rect -2189 -49440 1651 -45600
rect -2189 -53760 1651 -49920
<< metal5 >>
rect -429 53784 -109 54000
rect 2011 53839 2331 54000
rect -2213 53760 1675 53784
rect -2213 49920 -2189 53760
rect 1651 49920 1675 53760
rect -2213 49896 1675 49920
rect -429 49464 -109 49896
rect 2011 49841 2053 53839
rect 2289 49841 2331 53839
rect 2011 49519 2331 49841
rect -2213 49440 1675 49464
rect -2213 45600 -2189 49440
rect 1651 45600 1675 49440
rect -2213 45576 1675 45600
rect -429 45144 -109 45576
rect 2011 45521 2053 49519
rect 2289 45521 2331 49519
rect 2011 45199 2331 45521
rect -2213 45120 1675 45144
rect -2213 41280 -2189 45120
rect 1651 41280 1675 45120
rect -2213 41256 1675 41280
rect -429 40824 -109 41256
rect 2011 41201 2053 45199
rect 2289 41201 2331 45199
rect 2011 40879 2331 41201
rect -2213 40800 1675 40824
rect -2213 36960 -2189 40800
rect 1651 36960 1675 40800
rect -2213 36936 1675 36960
rect -429 36504 -109 36936
rect 2011 36881 2053 40879
rect 2289 36881 2331 40879
rect 2011 36559 2331 36881
rect -2213 36480 1675 36504
rect -2213 32640 -2189 36480
rect 1651 32640 1675 36480
rect -2213 32616 1675 32640
rect -429 32184 -109 32616
rect 2011 32561 2053 36559
rect 2289 32561 2331 36559
rect 2011 32239 2331 32561
rect -2213 32160 1675 32184
rect -2213 28320 -2189 32160
rect 1651 28320 1675 32160
rect -2213 28296 1675 28320
rect -429 27864 -109 28296
rect 2011 28241 2053 32239
rect 2289 28241 2331 32239
rect 2011 27919 2331 28241
rect -2213 27840 1675 27864
rect -2213 24000 -2189 27840
rect 1651 24000 1675 27840
rect -2213 23976 1675 24000
rect -429 23544 -109 23976
rect 2011 23921 2053 27919
rect 2289 23921 2331 27919
rect 2011 23599 2331 23921
rect -2213 23520 1675 23544
rect -2213 19680 -2189 23520
rect 1651 19680 1675 23520
rect -2213 19656 1675 19680
rect -429 19224 -109 19656
rect 2011 19601 2053 23599
rect 2289 19601 2331 23599
rect 2011 19279 2331 19601
rect -2213 19200 1675 19224
rect -2213 15360 -2189 19200
rect 1651 15360 1675 19200
rect -2213 15336 1675 15360
rect -429 14904 -109 15336
rect 2011 15281 2053 19279
rect 2289 15281 2331 19279
rect 2011 14959 2331 15281
rect -2213 14880 1675 14904
rect -2213 11040 -2189 14880
rect 1651 11040 1675 14880
rect -2213 11016 1675 11040
rect -429 10584 -109 11016
rect 2011 10961 2053 14959
rect 2289 10961 2331 14959
rect 2011 10639 2331 10961
rect -2213 10560 1675 10584
rect -2213 6720 -2189 10560
rect 1651 6720 1675 10560
rect -2213 6696 1675 6720
rect -429 6264 -109 6696
rect 2011 6641 2053 10639
rect 2289 6641 2331 10639
rect 2011 6319 2331 6641
rect -2213 6240 1675 6264
rect -2213 2400 -2189 6240
rect 1651 2400 1675 6240
rect -2213 2376 1675 2400
rect -429 1944 -109 2376
rect 2011 2321 2053 6319
rect 2289 2321 2331 6319
rect 2011 1999 2331 2321
rect -2213 1920 1675 1944
rect -2213 -1920 -2189 1920
rect 1651 -1920 1675 1920
rect -2213 -1944 1675 -1920
rect -429 -2376 -109 -1944
rect 2011 -1999 2053 1999
rect 2289 -1999 2331 1999
rect 2011 -2321 2331 -1999
rect -2213 -2400 1675 -2376
rect -2213 -6240 -2189 -2400
rect 1651 -6240 1675 -2400
rect -2213 -6264 1675 -6240
rect -429 -6696 -109 -6264
rect 2011 -6319 2053 -2321
rect 2289 -6319 2331 -2321
rect 2011 -6641 2331 -6319
rect -2213 -6720 1675 -6696
rect -2213 -10560 -2189 -6720
rect 1651 -10560 1675 -6720
rect -2213 -10584 1675 -10560
rect -429 -11016 -109 -10584
rect 2011 -10639 2053 -6641
rect 2289 -10639 2331 -6641
rect 2011 -10961 2331 -10639
rect -2213 -11040 1675 -11016
rect -2213 -14880 -2189 -11040
rect 1651 -14880 1675 -11040
rect -2213 -14904 1675 -14880
rect -429 -15336 -109 -14904
rect 2011 -14959 2053 -10961
rect 2289 -14959 2331 -10961
rect 2011 -15281 2331 -14959
rect -2213 -15360 1675 -15336
rect -2213 -19200 -2189 -15360
rect 1651 -19200 1675 -15360
rect -2213 -19224 1675 -19200
rect -429 -19656 -109 -19224
rect 2011 -19279 2053 -15281
rect 2289 -19279 2331 -15281
rect 2011 -19601 2331 -19279
rect -2213 -19680 1675 -19656
rect -2213 -23520 -2189 -19680
rect 1651 -23520 1675 -19680
rect -2213 -23544 1675 -23520
rect -429 -23976 -109 -23544
rect 2011 -23599 2053 -19601
rect 2289 -23599 2331 -19601
rect 2011 -23921 2331 -23599
rect -2213 -24000 1675 -23976
rect -2213 -27840 -2189 -24000
rect 1651 -27840 1675 -24000
rect -2213 -27864 1675 -27840
rect -429 -28296 -109 -27864
rect 2011 -27919 2053 -23921
rect 2289 -27919 2331 -23921
rect 2011 -28241 2331 -27919
rect -2213 -28320 1675 -28296
rect -2213 -32160 -2189 -28320
rect 1651 -32160 1675 -28320
rect -2213 -32184 1675 -32160
rect -429 -32616 -109 -32184
rect 2011 -32239 2053 -28241
rect 2289 -32239 2331 -28241
rect 2011 -32561 2331 -32239
rect -2213 -32640 1675 -32616
rect -2213 -36480 -2189 -32640
rect 1651 -36480 1675 -32640
rect -2213 -36504 1675 -36480
rect -429 -36936 -109 -36504
rect 2011 -36559 2053 -32561
rect 2289 -36559 2331 -32561
rect 2011 -36881 2331 -36559
rect -2213 -36960 1675 -36936
rect -2213 -40800 -2189 -36960
rect 1651 -40800 1675 -36960
rect -2213 -40824 1675 -40800
rect -429 -41256 -109 -40824
rect 2011 -40879 2053 -36881
rect 2289 -40879 2331 -36881
rect 2011 -41201 2331 -40879
rect -2213 -41280 1675 -41256
rect -2213 -45120 -2189 -41280
rect 1651 -45120 1675 -41280
rect -2213 -45144 1675 -45120
rect -429 -45576 -109 -45144
rect 2011 -45199 2053 -41201
rect 2289 -45199 2331 -41201
rect 2011 -45521 2331 -45199
rect -2213 -45600 1675 -45576
rect -2213 -49440 -2189 -45600
rect 1651 -49440 1675 -45600
rect -2213 -49464 1675 -49440
rect -429 -49896 -109 -49464
rect 2011 -49519 2053 -45521
rect 2289 -49519 2331 -45521
rect 2011 -49841 2331 -49519
rect -2213 -49920 1675 -49896
rect -2213 -53760 -2189 -49920
rect 1651 -53760 1675 -49920
rect -2213 -53784 1675 -53760
rect -429 -54000 -109 -53784
rect 2011 -53839 2053 -49841
rect 2289 -53839 2331 -49841
rect 2011 -54000 2331 -53839
<< properties >>
string FIXED_BBOX -2309 49800 1771 53880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 19.6 l 19.6 val 783.216 carea 2.00 cperi 0.19 nx 1 ny 25 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
