magic
tech sky130A
magscale 1 2
timestamp 1645495691
<< error_p >>
rect 2634 -36612 2930 36612
rect 2954 30781 3250 36563
rect 2954 30559 3274 30781
rect 2954 30239 3274 30461
rect 2954 24679 3250 30239
rect 2954 24457 3274 24679
rect 2954 24137 3274 24359
rect 2954 18577 3250 24137
rect 2954 18355 3274 18577
rect 2954 18035 3274 18257
rect 2954 12475 3250 18035
rect 2954 12253 3274 12475
rect 2954 11933 3274 12155
rect 2954 6373 3250 11933
rect 2954 6151 3274 6373
rect 2954 5831 3274 6053
rect 2954 271 3250 5831
rect 2954 49 3274 271
rect 2954 -271 3274 -49
rect 2954 -5831 3250 -271
rect 2954 -6053 3274 -5831
rect 2954 -6373 3274 -6151
rect 2954 -11933 3250 -6373
rect 2954 -12155 3274 -11933
rect 2954 -12475 3274 -12253
rect 2954 -18035 3250 -12475
rect 2954 -18257 3274 -18035
rect 2954 -18577 3274 -18355
rect 2954 -24137 3250 -18577
rect 2954 -24359 3274 -24137
rect 2954 -24679 3274 -24457
rect 2954 -30239 3250 -24679
rect 2954 -30461 3274 -30239
rect 2954 -30781 3274 -30559
rect 2954 -36563 3250 -30781
<< metal4 >>
rect -3252 36521 3252 36562
rect -3252 30601 2996 36521
rect 3232 30601 3252 36521
rect -3252 30560 3252 30601
rect -3252 30419 3252 30460
rect -3252 24499 2996 30419
rect 3232 24499 3252 30419
rect -3252 24458 3252 24499
rect -3252 24317 3252 24358
rect -3252 18397 2996 24317
rect 3232 18397 3252 24317
rect -3252 18356 3252 18397
rect -3252 18215 3252 18256
rect -3252 12295 2996 18215
rect 3232 12295 3252 18215
rect -3252 12254 3252 12295
rect -3252 12113 3252 12154
rect -3252 6193 2996 12113
rect 3232 6193 3252 12113
rect -3252 6152 3252 6193
rect -3252 6011 3252 6052
rect -3252 91 2996 6011
rect 3232 91 3252 6011
rect -3252 50 3252 91
rect -3252 -91 3252 -50
rect -3252 -6011 2996 -91
rect 3232 -6011 3252 -91
rect -3252 -6052 3252 -6011
rect -3252 -6193 3252 -6152
rect -3252 -12113 2996 -6193
rect 3232 -12113 3252 -6193
rect -3252 -12154 3252 -12113
rect -3252 -12295 3252 -12254
rect -3252 -18215 2996 -12295
rect 3232 -18215 3252 -12295
rect -3252 -18256 3252 -18215
rect -3252 -18397 3252 -18356
rect -3252 -24317 2996 -18397
rect 3232 -24317 3252 -18397
rect -3252 -24358 3252 -24317
rect -3252 -24499 3252 -24458
rect -3252 -30419 2996 -24499
rect 3232 -30419 3252 -24499
rect -3252 -30460 3252 -30419
rect -3252 -30601 3252 -30560
rect -3252 -36521 2996 -30601
rect 3232 -36521 3252 -30601
rect -3252 -36562 3252 -36521
<< via4 >>
rect 2996 30601 3232 36521
rect 2996 24499 3232 30419
rect 2996 18397 3232 24317
rect 2996 12295 3232 18215
rect 2996 6193 3232 12113
rect 2996 91 3232 6011
rect 2996 -6011 3232 -91
rect 2996 -12113 3232 -6193
rect 2996 -18215 3232 -12295
rect 2996 -24317 3232 -18397
rect 2996 -30419 3232 -24499
rect 2996 -36521 3232 -30601
<< mimcap2 >>
rect -3152 36422 2650 36462
rect -3152 30700 -3112 36422
rect 2610 30700 2650 36422
rect -3152 30660 2650 30700
rect -3152 30320 2650 30360
rect -3152 24598 -3112 30320
rect 2610 24598 2650 30320
rect -3152 24558 2650 24598
rect -3152 24218 2650 24258
rect -3152 18496 -3112 24218
rect 2610 18496 2650 24218
rect -3152 18456 2650 18496
rect -3152 18116 2650 18156
rect -3152 12394 -3112 18116
rect 2610 12394 2650 18116
rect -3152 12354 2650 12394
rect -3152 12014 2650 12054
rect -3152 6292 -3112 12014
rect 2610 6292 2650 12014
rect -3152 6252 2650 6292
rect -3152 5912 2650 5952
rect -3152 190 -3112 5912
rect 2610 190 2650 5912
rect -3152 150 2650 190
rect -3152 -190 2650 -150
rect -3152 -5912 -3112 -190
rect 2610 -5912 2650 -190
rect -3152 -5952 2650 -5912
rect -3152 -6292 2650 -6252
rect -3152 -12014 -3112 -6292
rect 2610 -12014 2650 -6292
rect -3152 -12054 2650 -12014
rect -3152 -12394 2650 -12354
rect -3152 -18116 -3112 -12394
rect 2610 -18116 2650 -12394
rect -3152 -18156 2650 -18116
rect -3152 -18496 2650 -18456
rect -3152 -24218 -3112 -18496
rect 2610 -24218 2650 -18496
rect -3152 -24258 2650 -24218
rect -3152 -24598 2650 -24558
rect -3152 -30320 -3112 -24598
rect 2610 -30320 2650 -24598
rect -3152 -30360 2650 -30320
rect -3152 -30700 2650 -30660
rect -3152 -36422 -3112 -30700
rect 2610 -36422 2650 -30700
rect -3152 -36462 2650 -36422
<< mimcap2contact >>
rect -3112 30700 2610 36422
rect -3112 24598 2610 30320
rect -3112 18496 2610 24218
rect -3112 12394 2610 18116
rect -3112 6292 2610 12014
rect -3112 190 2610 5912
rect -3112 -5912 2610 -190
rect -3112 -12014 2610 -6292
rect -3112 -18116 2610 -12394
rect -3112 -24218 2610 -18496
rect -3112 -30320 2610 -24598
rect -3112 -36422 2610 -30700
<< metal5 >>
rect -411 36446 -91 36612
rect 2610 36446 2930 36612
rect -3136 36422 2930 36446
rect -3136 30700 -3112 36422
rect 2610 30700 2930 36422
rect -3136 30676 2930 30700
rect -411 30344 -91 30676
rect 2610 30344 2930 30676
rect 2954 36521 3274 36563
rect 2954 30601 2996 36521
rect 3232 30601 3274 36521
rect 2954 30559 3274 30601
rect -3136 30320 2930 30344
rect -3136 24598 -3112 30320
rect 2610 24598 2930 30320
rect -3136 24574 2930 24598
rect -411 24242 -91 24574
rect 2610 24242 2930 24574
rect 2954 30419 3274 30461
rect 2954 24499 2996 30419
rect 3232 24499 3274 30419
rect 2954 24457 3274 24499
rect -3136 24218 2930 24242
rect -3136 18496 -3112 24218
rect 2610 18496 2930 24218
rect -3136 18472 2930 18496
rect -411 18140 -91 18472
rect 2610 18140 2930 18472
rect 2954 24317 3274 24359
rect 2954 18397 2996 24317
rect 3232 18397 3274 24317
rect 2954 18355 3274 18397
rect -3136 18116 2930 18140
rect -3136 12394 -3112 18116
rect 2610 12394 2930 18116
rect -3136 12370 2930 12394
rect -411 12038 -91 12370
rect 2610 12038 2930 12370
rect 2954 18215 3274 18257
rect 2954 12295 2996 18215
rect 3232 12295 3274 18215
rect 2954 12253 3274 12295
rect -3136 12014 2930 12038
rect -3136 6292 -3112 12014
rect 2610 6292 2930 12014
rect -3136 6268 2930 6292
rect -411 5936 -91 6268
rect 2610 5936 2930 6268
rect 2954 12113 3274 12155
rect 2954 6193 2996 12113
rect 3232 6193 3274 12113
rect 2954 6151 3274 6193
rect -3136 5912 2930 5936
rect -3136 190 -3112 5912
rect 2610 190 2930 5912
rect -3136 166 2930 190
rect -411 -166 -91 166
rect 2610 -166 2930 166
rect 2954 6011 3274 6053
rect 2954 91 2996 6011
rect 3232 91 3274 6011
rect 2954 49 3274 91
rect -3136 -190 2930 -166
rect -3136 -5912 -3112 -190
rect 2610 -5912 2930 -190
rect -3136 -5936 2930 -5912
rect -411 -6268 -91 -5936
rect 2610 -6268 2930 -5936
rect 2954 -91 3274 -49
rect 2954 -6011 2996 -91
rect 3232 -6011 3274 -91
rect 2954 -6053 3274 -6011
rect -3136 -6292 2930 -6268
rect -3136 -12014 -3112 -6292
rect 2610 -12014 2930 -6292
rect -3136 -12038 2930 -12014
rect -411 -12370 -91 -12038
rect 2610 -12370 2930 -12038
rect 2954 -6193 3274 -6151
rect 2954 -12113 2996 -6193
rect 3232 -12113 3274 -6193
rect 2954 -12155 3274 -12113
rect -3136 -12394 2930 -12370
rect -3136 -18116 -3112 -12394
rect 2610 -18116 2930 -12394
rect -3136 -18140 2930 -18116
rect -411 -18472 -91 -18140
rect 2610 -18472 2930 -18140
rect 2954 -12295 3274 -12253
rect 2954 -18215 2996 -12295
rect 3232 -18215 3274 -12295
rect 2954 -18257 3274 -18215
rect -3136 -18496 2930 -18472
rect -3136 -24218 -3112 -18496
rect 2610 -24218 2930 -18496
rect -3136 -24242 2930 -24218
rect -411 -24574 -91 -24242
rect 2610 -24574 2930 -24242
rect 2954 -18397 3274 -18355
rect 2954 -24317 2996 -18397
rect 3232 -24317 3274 -18397
rect 2954 -24359 3274 -24317
rect -3136 -24598 2930 -24574
rect -3136 -30320 -3112 -24598
rect 2610 -30320 2930 -24598
rect -3136 -30344 2930 -30320
rect -411 -30676 -91 -30344
rect 2610 -30676 2930 -30344
rect 2954 -24499 3274 -24457
rect 2954 -30419 2996 -24499
rect 3232 -30419 3274 -24499
rect 2954 -30461 3274 -30419
rect -3136 -30700 2930 -30676
rect -3136 -36422 -3112 -30700
rect 2610 -36422 2930 -30700
rect -3136 -36446 2930 -36422
rect -411 -36612 -91 -36446
rect 2610 -36612 2930 -36446
rect 2954 -30601 3274 -30559
rect 2954 -36521 2996 -30601
rect 3232 -36521 3274 -30601
rect 2954 -36563 3274 -36521
<< properties >>
string FIXED_BBOX -3252 30560 2750 36562
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 29.008 l 29.008 val 1.704k carea 2.00 cperi 0.19 nx 1 ny 12 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
