magic
tech sky130A
magscale 1 2
timestamp 1655563127
<< nwell >>
rect -683 -1019 683 1019
<< pmos >>
rect -487 -800 -287 800
rect -229 -800 -29 800
rect 29 -800 229 800
rect 287 -800 487 800
<< pdiff >>
rect -545 788 -487 800
rect -545 -788 -533 788
rect -499 -788 -487 788
rect -545 -800 -487 -788
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
rect 487 788 545 800
rect 487 -788 499 788
rect 533 -788 545 788
rect 487 -800 545 -788
<< pdiffc >>
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
<< nsubdiff >>
rect -647 949 -551 983
rect 551 949 647 983
rect -647 887 -613 949
rect 613 887 647 949
rect -647 -949 -613 -887
rect 613 -949 647 -887
rect -647 -983 -551 -949
rect 551 -983 647 -949
<< nsubdiffcont >>
rect -551 949 551 983
rect -647 -887 -613 887
rect 613 -887 647 887
rect -551 -983 551 -949
<< poly >>
rect -487 881 -287 897
rect -487 847 -471 881
rect -303 847 -287 881
rect -487 800 -287 847
rect -229 881 -29 897
rect -229 847 -213 881
rect -45 847 -29 881
rect -229 800 -29 847
rect 29 881 229 897
rect 29 847 45 881
rect 213 847 229 881
rect 29 800 229 847
rect 287 881 487 897
rect 287 847 303 881
rect 471 847 487 881
rect 287 800 487 847
rect -487 -847 -287 -800
rect -487 -881 -471 -847
rect -303 -881 -287 -847
rect -487 -897 -287 -881
rect -229 -847 -29 -800
rect -229 -881 -213 -847
rect -45 -881 -29 -847
rect -229 -897 -29 -881
rect 29 -847 229 -800
rect 29 -881 45 -847
rect 213 -881 229 -847
rect 29 -897 229 -881
rect 287 -847 487 -800
rect 287 -881 303 -847
rect 471 -881 487 -847
rect 287 -897 487 -881
<< polycont >>
rect -471 847 -303 881
rect -213 847 -45 881
rect 45 847 213 881
rect 303 847 471 881
rect -471 -881 -303 -847
rect -213 -881 -45 -847
rect 45 -881 213 -847
rect 303 -881 471 -847
<< locali >>
rect -647 949 -551 983
rect 551 949 647 983
rect -647 887 -613 949
rect 613 887 647 949
rect -487 847 -471 881
rect -303 847 -287 881
rect -229 847 -213 881
rect -45 847 -29 881
rect 29 847 45 881
rect 213 847 229 881
rect 287 847 303 881
rect 471 847 487 881
rect -533 788 -499 804
rect -533 -804 -499 -788
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
rect 499 788 533 804
rect 499 -804 533 -788
rect -487 -881 -471 -847
rect -303 -881 -287 -847
rect -229 -881 -213 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 213 -881 229 -847
rect 287 -881 303 -847
rect 471 -881 487 -847
rect -647 -949 -613 -887
rect 613 -949 647 -887
rect -647 -983 -551 -949
rect 551 -983 647 -949
<< viali >>
rect -471 847 -303 881
rect -213 847 -45 881
rect 45 847 213 881
rect 303 847 471 881
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
rect -471 -881 -303 -847
rect -213 -881 -45 -847
rect 45 -881 213 -847
rect 303 -881 471 -847
<< metal1 >>
rect -483 881 -291 887
rect -483 847 -471 881
rect -303 847 -291 881
rect -483 841 -291 847
rect -225 881 -33 887
rect -225 847 -213 881
rect -45 847 -33 881
rect -225 841 -33 847
rect 33 881 225 887
rect 33 847 45 881
rect 213 847 225 881
rect 33 841 225 847
rect 291 881 483 887
rect 291 847 303 881
rect 471 847 483 881
rect 291 841 483 847
rect -539 788 -493 800
rect -539 -788 -533 788
rect -499 -788 -493 788
rect -539 -800 -493 -788
rect -281 788 -235 800
rect -281 -788 -275 788
rect -241 -788 -235 788
rect -281 -800 -235 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 235 788 281 800
rect 235 -788 241 788
rect 275 -788 281 788
rect 235 -800 281 -788
rect 493 788 539 800
rect 493 -788 499 788
rect 533 -788 539 788
rect 493 -800 539 -788
rect -483 -847 -291 -841
rect -483 -881 -471 -847
rect -303 -881 -291 -847
rect -483 -887 -291 -881
rect -225 -847 -33 -841
rect -225 -881 -213 -847
rect -45 -881 -33 -847
rect -225 -887 -33 -881
rect 33 -847 225 -841
rect 33 -881 45 -847
rect 213 -881 225 -847
rect 33 -887 225 -881
rect 291 -847 483 -841
rect 291 -881 303 -847
rect 471 -881 483 -847
rect 291 -887 483 -881
<< properties >>
string FIXED_BBOX -630 -966 630 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
