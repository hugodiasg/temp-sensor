magic
tech sky130A
magscale 1 2
timestamp 1661301161
<< nwell >>
rect -812 -319 812 319
<< pmos >>
rect -616 -100 -416 100
rect -358 -100 -158 100
rect -100 -100 100 100
rect 158 -100 358 100
rect 416 -100 616 100
<< pdiff >>
rect -674 88 -616 100
rect -674 -88 -662 88
rect -628 -88 -616 88
rect -674 -100 -616 -88
rect -416 88 -358 100
rect -416 -88 -404 88
rect -370 -88 -358 88
rect -416 -100 -358 -88
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
rect 358 88 416 100
rect 358 -88 370 88
rect 404 -88 416 88
rect 358 -100 416 -88
rect 616 88 674 100
rect 616 -88 628 88
rect 662 -88 674 88
rect 616 -100 674 -88
<< pdiffc >>
rect -662 -88 -628 88
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
rect 628 -88 662 88
<< nsubdiff >>
rect -776 249 -680 283
rect 680 249 776 283
rect -776 187 -742 249
rect 742 187 776 249
rect -776 -249 -742 -187
rect 742 -249 776 -187
rect -776 -283 -680 -249
rect 680 -283 776 -249
<< nsubdiffcont >>
rect -680 249 680 283
rect -776 -187 -742 187
rect 742 -187 776 187
rect -680 -283 680 -249
<< poly >>
rect -616 181 -416 197
rect -616 147 -600 181
rect -432 147 -416 181
rect -616 100 -416 147
rect -358 181 -158 197
rect -358 147 -342 181
rect -174 147 -158 181
rect -358 100 -158 147
rect -100 181 100 197
rect -100 147 -84 181
rect 84 147 100 181
rect -100 100 100 147
rect 158 181 358 197
rect 158 147 174 181
rect 342 147 358 181
rect 158 100 358 147
rect 416 181 616 197
rect 416 147 432 181
rect 600 147 616 181
rect 416 100 616 147
rect -616 -147 -416 -100
rect -616 -181 -600 -147
rect -432 -181 -416 -147
rect -616 -197 -416 -181
rect -358 -147 -158 -100
rect -358 -181 -342 -147
rect -174 -181 -158 -147
rect -358 -197 -158 -181
rect -100 -147 100 -100
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -100 -197 100 -181
rect 158 -147 358 -100
rect 158 -181 174 -147
rect 342 -181 358 -147
rect 158 -197 358 -181
rect 416 -147 616 -100
rect 416 -181 432 -147
rect 600 -181 616 -147
rect 416 -197 616 -181
<< polycont >>
rect -600 147 -432 181
rect -342 147 -174 181
rect -84 147 84 181
rect 174 147 342 181
rect 432 147 600 181
rect -600 -181 -432 -147
rect -342 -181 -174 -147
rect -84 -181 84 -147
rect 174 -181 342 -147
rect 432 -181 600 -147
<< locali >>
rect -776 249 -680 283
rect 680 249 776 283
rect 742 187 776 249
rect -616 147 -600 181
rect -432 147 -416 181
rect -358 147 -342 181
rect -174 147 -158 181
rect -100 147 -84 181
rect 84 147 100 181
rect 158 147 174 181
rect 342 147 358 181
rect 416 147 432 181
rect 600 147 616 181
rect -662 88 -628 104
rect -662 -104 -628 -88
rect -404 88 -370 104
rect -404 -104 -370 -88
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect 370 88 404 104
rect 370 -104 404 -88
rect 628 88 662 104
rect 628 -104 662 -88
rect -616 -181 -600 -147
rect -432 -181 -416 -147
rect -358 -181 -342 -147
rect -174 -181 -158 -147
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect 158 -181 174 -147
rect 342 -181 358 -147
rect 416 -181 432 -147
rect 600 -181 616 -147
rect 742 -249 776 -187
rect -776 -283 -680 -249
rect 680 -283 776 -249
<< viali >>
rect -776 187 -742 249
rect -776 -187 -742 187
rect -600 147 -432 181
rect -342 147 -174 181
rect -84 147 84 181
rect 174 147 342 181
rect 432 147 600 181
rect -662 1 -628 71
rect -404 -35 -370 35
rect -146 1 -112 71
rect 112 -35 146 35
rect 370 1 404 71
rect 628 -35 662 35
rect -600 -181 -432 -147
rect -342 -181 -174 -147
rect -84 -181 84 -147
rect 174 -181 342 -147
rect 432 -181 600 -147
rect -776 -249 -742 -187
<< metal1 >>
rect -782 249 -736 261
rect -782 -249 -776 249
rect -742 -249 -736 249
rect -612 181 -420 187
rect -612 147 -600 181
rect -432 147 -420 181
rect -612 141 -420 147
rect -354 181 -162 187
rect -354 147 -342 181
rect -174 147 -162 181
rect -354 141 -162 147
rect -96 181 96 187
rect -96 147 -84 181
rect 84 147 96 181
rect -96 141 96 147
rect 162 181 354 187
rect 162 147 174 181
rect 342 147 354 181
rect 162 141 354 147
rect 420 181 612 187
rect 420 147 432 181
rect 600 147 612 181
rect 420 141 612 147
rect -668 71 -622 83
rect -668 1 -662 71
rect -628 1 -622 71
rect -152 71 -106 83
rect -668 -11 -622 1
rect -410 35 -364 47
rect -410 -35 -404 35
rect -370 -35 -364 35
rect -152 1 -146 71
rect -112 1 -106 71
rect 364 71 410 83
rect -152 -11 -106 1
rect 106 35 152 47
rect -410 -47 -364 -35
rect 106 -35 112 35
rect 146 -35 152 35
rect 364 1 370 71
rect 404 1 410 71
rect 364 -11 410 1
rect 622 35 668 47
rect 106 -47 152 -35
rect 622 -35 628 35
rect 662 -35 668 35
rect 622 -47 668 -35
rect -612 -147 -420 -141
rect -612 -181 -600 -147
rect -432 -181 -420 -147
rect -612 -187 -420 -181
rect -354 -147 -162 -141
rect -354 -181 -342 -147
rect -174 -181 -162 -147
rect -354 -187 -162 -181
rect -96 -147 96 -141
rect -96 -181 -84 -147
rect 84 -181 96 -147
rect -96 -187 96 -181
rect 162 -147 354 -141
rect 162 -181 174 -147
rect 342 -181 354 -147
rect 162 -187 354 -181
rect 420 -147 612 -141
rect 420 -181 432 -147
rect 600 -181 612 -147
rect 420 -187 612 -181
rect -782 -261 -736 -249
<< properties >>
string FIXED_BBOX -759 -266 759 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 100 viagt 0
<< end >>
