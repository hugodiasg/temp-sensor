** sch_path: /foss/designs/temp-sensor/sigma-delta_modulator/xschem/sigma_tb-tran.sch
**.subckt sigma_tb-tran
vin in1 GND 1.2
vpwr vpwr GND 1.8
V3 clk GND pulse 0 1.8 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 '
vd vd GND 1.8
vin1 in2 GND 1.3
vin2 in3 GND 1.4
Bvts in_linear GND v=200*time+1.2
XC1 net1 net2 sky130_fd_pr__cap_mim_m3_1 W=27.196 L=27.196 MF=1 m=1
x1 vpwr clk out1 in1 vpwr GND vd sigma-delta
x2 vpwr clk out2 in2 vpwr GND vd sigma-delta
x3 vpwr clk out3 in3 vpwr GND vd sigma-delta
**** begin user architecture code

*cmd step stop
*PULSE ( V1 V2 TD TR TF PW PER PHASE)
.control
destroy all
save all
set color0=white
set color1=black
tran 10n 10u
*tran 10n 1m
run

*plot in_linear out1
plot in1 out1
plot in2 out2
plot in3 out3

.endc

 .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sym # of
*+ pins=7
** sym_path: /foss/designs/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sym
** sch_path: /foss/designs/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sch
.subckt sigma-delta vpwr clk out in reset_b_dff gnd vd
*.ipin in
*.iopin gnd
*.iopin clk
*.iopin out
*.iopin reset_b_dff
*.iopin vpwr
*.iopin vd
XR2 Q in_int gnd sky130_fd_pr__res_xhigh_po_0p35 L=36 mult=1 m=1
XR1 in_int in gnd sky130_fd_pr__res_xhigh_po_0p35 L=36 mult=1 m=1
XN1 out_comp in_comp gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XP1 out_comp in_comp vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x1 clk out_comp reset_b_dff GND GND VPWR VPWR Q out sky130_fd_sc_hd__dfrbp_1
XR3 in_comp in_int gnd sky130_fd_pr__res_xhigh_po_0p35 L=18 mult=1 m=1
**** begin user architecture code

.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


**** end user architecture code
XC1 in_int gnd sky130_fd_pr__cap_mim_m3_1 W=27.196 L=27.196 MF=1 m=1
XC2 in_comp gnd sky130_fd_pr__cap_mim_m3_1 W=27.196 L=27.196 MF=1 m=1
.ends

.GLOBAL GND
.end
