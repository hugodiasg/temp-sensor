magic
tech sky130A
magscale 1 2
timestamp 1700192422
<< nwell >>
rect 5647 5567 12813 6253
rect 207 3627 4233 5293
rect 167 2307 3393 3373
rect 14320 3050 14740 3060
rect 14320 2820 16752 3050
rect 14560 2729 16752 2820
rect 17014 2594 17436 3632
<< pwell >>
rect 5960 29220 6362 31416
rect 680 10340 1102 11160
rect 5700 4680 12092 5300
rect 5780 3840 12560 4460
rect 15501 2625 15687 2669
rect 16231 2625 16702 2671
rect 14599 2489 16702 2625
rect 14627 2451 14661 2489
rect 0 160 3392 2080
rect 17014 1924 17436 2544
<< nmos >>
rect 876 10550 906 10950
rect 5884 4882 6084 5082
rect 6142 4882 6342 5082
rect 6400 4882 6600 5082
rect 6658 4882 6858 5082
rect 6916 4882 7116 5082
rect 7174 4882 7374 5082
rect 7432 4882 7632 5082
rect 7690 4882 7890 5082
rect 7948 4882 8148 5082
rect 8206 4882 8406 5082
rect 8464 4882 8664 5082
rect 8722 4882 8922 5082
rect 8980 4882 9180 5082
rect 9238 4882 9438 5082
rect 9496 4882 9696 5082
rect 9754 4882 9954 5082
rect 10012 4882 10212 5082
rect 10270 4882 10470 5082
rect 10528 4882 10728 5082
rect 10786 4882 10986 5082
rect 11044 4882 11244 5082
rect 11302 4882 11502 5082
rect 5978 4048 6178 4248
rect 6236 4048 6436 4248
rect 6494 4048 6694 4248
rect 6898 4048 7098 4248
rect 7156 4048 7356 4248
rect 7414 4048 7614 4248
rect 7672 4048 7872 4248
rect 7930 4048 8130 4248
rect 8188 4048 8388 4248
rect 8446 4048 8646 4248
rect 8704 4048 8904 4248
rect 8962 4048 9162 4248
rect 9220 4048 9420 4248
rect 9478 4048 9678 4248
rect 9736 4048 9936 4248
rect 9994 4048 10194 4248
rect 10252 4048 10452 4248
rect 10510 4048 10710 4248
rect 10768 4048 10968 4248
rect 11026 4048 11226 4248
rect 11284 4048 11484 4248
rect 11542 4048 11742 4248
rect 11800 4048 12000 4248
rect 12058 4048 12258 4248
rect 17210 2134 17240 2334
rect 218 1672 418 1872
rect 598 1672 798 1872
rect 978 1672 1178 1872
rect 1358 1672 1558 1872
rect 1738 1672 1938 1872
rect 2118 1672 2318 1872
rect 2498 1672 2698 1872
rect 2878 1672 3078 1872
rect 218 1254 418 1454
rect 598 1254 798 1454
rect 978 1254 1178 1454
rect 1358 1254 1558 1454
rect 1738 1254 1938 1454
rect 2118 1254 2318 1454
rect 2498 1254 2698 1454
rect 2878 1254 3078 1454
rect 218 836 418 1036
rect 598 836 798 1036
rect 978 836 1178 1036
rect 1358 836 1558 1036
rect 1738 836 1938 1036
rect 2118 836 2318 1036
rect 2498 836 2698 1036
rect 2878 836 3078 1036
rect 218 418 418 618
rect 598 418 798 618
rect 978 418 1178 618
rect 1358 418 1558 618
rect 1738 418 1938 618
rect 2118 418 2318 618
rect 2498 418 2698 618
rect 2878 418 3078 618
<< scnmos >>
rect 14677 2515 14707 2599
rect 14761 2515 14791 2599
rect 15016 2515 15046 2599
rect 15111 2515 15141 2587
rect 15207 2515 15237 2587
rect 15373 2515 15403 2599
rect 15445 2515 15475 2599
rect 15577 2515 15607 2643
rect 15676 2515 15706 2587
rect 15785 2515 15815 2587
rect 15881 2515 15911 2599
rect 16030 2515 16060 2599
rect 16121 2515 16151 2599
rect 16309 2515 16339 2645
rect 16497 2515 16527 2599
rect 16594 2515 16624 2645
<< pmos >>
rect 5854 5800 6054 6000
rect 6112 5800 6312 6000
rect 6370 5800 6570 6000
rect 6628 5800 6828 6000
rect 6886 5800 7086 6000
rect 7144 5800 7344 6000
rect 7514 5800 7714 6000
rect 7894 5800 8094 6000
rect 8152 5800 8352 6000
rect 8410 5800 8610 6000
rect 8668 5800 8868 6000
rect 8926 5800 9126 6000
rect 9314 5800 9514 6000
rect 9572 5800 9772 6000
rect 9830 5800 10030 6000
rect 10088 5800 10288 6000
rect 10346 5800 10546 6000
rect 10734 5800 10934 6000
rect 11114 5800 11314 6000
rect 11372 5800 11572 6000
rect 11630 5800 11830 6000
rect 11888 5800 12088 6000
rect 12146 5800 12346 6000
rect 12404 5800 12604 6000
rect 1814 4580 2014 4980
rect 2194 4580 2394 4980
rect 2574 4580 3574 4980
rect 3754 4580 3954 4980
rect 434 3900 634 4300
rect 814 3900 1014 4300
rect 1072 3900 1272 4300
rect 1454 3900 1654 4300
rect 1712 3900 1912 4300
rect 1970 3900 2170 4300
rect 2228 3900 2428 4300
rect 2614 3900 2814 4300
rect 2872 3900 3072 4300
rect 3130 3900 3330 4300
rect 3388 3900 3588 4300
rect 3774 3900 3974 4300
rect 414 2660 614 3060
rect 794 2660 994 3060
rect 1052 2660 1252 3060
rect 1310 2660 1510 3060
rect 1568 2660 1768 3060
rect 1826 2660 2026 3060
rect 2084 2660 2284 3060
rect 2342 2660 2542 3060
rect 2600 2660 2800 3060
rect 2974 2660 3174 3060
rect 17210 2813 17240 3413
<< scpmoshvt >>
rect 14677 2831 14707 2959
rect 14761 2831 14791 2959
rect 15028 2881 15058 2965
rect 15120 2881 15150 2965
rect 15219 2881 15249 2965
rect 15359 2881 15389 2965
rect 15456 2881 15486 2965
rect 15653 2797 15683 2965
rect 15752 2881 15782 2965
rect 15838 2881 15868 2965
rect 15922 2881 15952 2965
rect 16030 2881 16060 2965
rect 16114 2881 16144 2965
rect 16278 2765 16308 2965
rect 16497 2837 16527 2965
rect 16594 2765 16624 2965
<< ndiff >>
rect 818 10938 876 10950
rect 818 10562 830 10938
rect 864 10562 876 10938
rect 818 10550 876 10562
rect 906 10938 964 10950
rect 906 10562 918 10938
rect 952 10562 964 10938
rect 906 10550 964 10562
rect 5826 5070 5884 5082
rect 5826 4894 5838 5070
rect 5872 4894 5884 5070
rect 5826 4882 5884 4894
rect 6084 5070 6142 5082
rect 6084 4894 6096 5070
rect 6130 4894 6142 5070
rect 6084 4882 6142 4894
rect 6342 5070 6400 5082
rect 6342 4894 6354 5070
rect 6388 4894 6400 5070
rect 6342 4882 6400 4894
rect 6600 5070 6658 5082
rect 6600 4894 6612 5070
rect 6646 4894 6658 5070
rect 6600 4882 6658 4894
rect 6858 5070 6916 5082
rect 6858 4894 6870 5070
rect 6904 4894 6916 5070
rect 6858 4882 6916 4894
rect 7116 5070 7174 5082
rect 7116 4894 7128 5070
rect 7162 4894 7174 5070
rect 7116 4882 7174 4894
rect 7374 5070 7432 5082
rect 7374 4894 7386 5070
rect 7420 4894 7432 5070
rect 7374 4882 7432 4894
rect 7632 5070 7690 5082
rect 7632 4894 7644 5070
rect 7678 4894 7690 5070
rect 7632 4882 7690 4894
rect 7890 5070 7948 5082
rect 7890 4894 7902 5070
rect 7936 4894 7948 5070
rect 7890 4882 7948 4894
rect 8148 5070 8206 5082
rect 8148 4894 8160 5070
rect 8194 4894 8206 5070
rect 8148 4882 8206 4894
rect 8406 5070 8464 5082
rect 8406 4894 8418 5070
rect 8452 4894 8464 5070
rect 8406 4882 8464 4894
rect 8664 5070 8722 5082
rect 8664 4894 8676 5070
rect 8710 4894 8722 5070
rect 8664 4882 8722 4894
rect 8922 5070 8980 5082
rect 8922 4894 8934 5070
rect 8968 4894 8980 5070
rect 8922 4882 8980 4894
rect 9180 5070 9238 5082
rect 9180 4894 9192 5070
rect 9226 4894 9238 5070
rect 9180 4882 9238 4894
rect 9438 5070 9496 5082
rect 9438 4894 9450 5070
rect 9484 4894 9496 5070
rect 9438 4882 9496 4894
rect 9696 5070 9754 5082
rect 9696 4894 9708 5070
rect 9742 4894 9754 5070
rect 9696 4882 9754 4894
rect 9954 5070 10012 5082
rect 9954 4894 9966 5070
rect 10000 4894 10012 5070
rect 9954 4882 10012 4894
rect 10212 5070 10270 5082
rect 10212 4894 10224 5070
rect 10258 4894 10270 5070
rect 10212 4882 10270 4894
rect 10470 5070 10528 5082
rect 10470 4894 10482 5070
rect 10516 4894 10528 5070
rect 10470 4882 10528 4894
rect 10728 5070 10786 5082
rect 10728 4894 10740 5070
rect 10774 4894 10786 5070
rect 10728 4882 10786 4894
rect 10986 5070 11044 5082
rect 10986 4894 10998 5070
rect 11032 4894 11044 5070
rect 10986 4882 11044 4894
rect 11244 5070 11302 5082
rect 11244 4894 11256 5070
rect 11290 4894 11302 5070
rect 11244 4882 11302 4894
rect 11502 5070 11560 5082
rect 11502 4894 11514 5070
rect 11548 4894 11560 5070
rect 11502 4882 11560 4894
rect 5920 4236 5978 4248
rect 5920 4060 5932 4236
rect 5966 4060 5978 4236
rect 5920 4048 5978 4060
rect 6178 4236 6236 4248
rect 6178 4060 6190 4236
rect 6224 4060 6236 4236
rect 6178 4048 6236 4060
rect 6436 4236 6494 4248
rect 6436 4060 6448 4236
rect 6482 4060 6494 4236
rect 6436 4048 6494 4060
rect 6694 4236 6752 4248
rect 6694 4060 6706 4236
rect 6740 4060 6752 4236
rect 6694 4048 6752 4060
rect 6840 4236 6898 4248
rect 6840 4060 6852 4236
rect 6886 4060 6898 4236
rect 6840 4048 6898 4060
rect 7098 4236 7156 4248
rect 7098 4060 7110 4236
rect 7144 4060 7156 4236
rect 7098 4048 7156 4060
rect 7356 4236 7414 4248
rect 7356 4060 7368 4236
rect 7402 4060 7414 4236
rect 7356 4048 7414 4060
rect 7614 4236 7672 4248
rect 7614 4060 7626 4236
rect 7660 4060 7672 4236
rect 7614 4048 7672 4060
rect 7872 4236 7930 4248
rect 7872 4060 7884 4236
rect 7918 4060 7930 4236
rect 7872 4048 7930 4060
rect 8130 4236 8188 4248
rect 8130 4060 8142 4236
rect 8176 4060 8188 4236
rect 8130 4048 8188 4060
rect 8388 4236 8446 4248
rect 8388 4060 8400 4236
rect 8434 4060 8446 4236
rect 8388 4048 8446 4060
rect 8646 4236 8704 4248
rect 8646 4060 8658 4236
rect 8692 4060 8704 4236
rect 8646 4048 8704 4060
rect 8904 4236 8962 4248
rect 8904 4060 8916 4236
rect 8950 4060 8962 4236
rect 8904 4048 8962 4060
rect 9162 4236 9220 4248
rect 9162 4060 9174 4236
rect 9208 4060 9220 4236
rect 9162 4048 9220 4060
rect 9420 4236 9478 4248
rect 9420 4060 9432 4236
rect 9466 4060 9478 4236
rect 9420 4048 9478 4060
rect 9678 4236 9736 4248
rect 9678 4060 9690 4236
rect 9724 4060 9736 4236
rect 9678 4048 9736 4060
rect 9936 4236 9994 4248
rect 9936 4060 9948 4236
rect 9982 4060 9994 4236
rect 9936 4048 9994 4060
rect 10194 4236 10252 4248
rect 10194 4060 10206 4236
rect 10240 4060 10252 4236
rect 10194 4048 10252 4060
rect 10452 4236 10510 4248
rect 10452 4060 10464 4236
rect 10498 4060 10510 4236
rect 10452 4048 10510 4060
rect 10710 4236 10768 4248
rect 10710 4060 10722 4236
rect 10756 4060 10768 4236
rect 10710 4048 10768 4060
rect 10968 4236 11026 4248
rect 10968 4060 10980 4236
rect 11014 4060 11026 4236
rect 10968 4048 11026 4060
rect 11226 4236 11284 4248
rect 11226 4060 11238 4236
rect 11272 4060 11284 4236
rect 11226 4048 11284 4060
rect 11484 4236 11542 4248
rect 11484 4060 11496 4236
rect 11530 4060 11542 4236
rect 11484 4048 11542 4060
rect 11742 4236 11800 4248
rect 11742 4060 11754 4236
rect 11788 4060 11800 4236
rect 11742 4048 11800 4060
rect 12000 4236 12058 4248
rect 12000 4060 12012 4236
rect 12046 4060 12058 4236
rect 12000 4048 12058 4060
rect 12258 4236 12316 4248
rect 12258 4060 12270 4236
rect 12304 4060 12316 4236
rect 12258 4048 12316 4060
rect 14625 2587 14677 2599
rect 14625 2553 14633 2587
rect 14667 2553 14677 2587
rect 14625 2515 14677 2553
rect 14707 2561 14761 2599
rect 14707 2527 14717 2561
rect 14751 2527 14761 2561
rect 14707 2515 14761 2527
rect 14791 2587 14843 2599
rect 14791 2553 14801 2587
rect 14835 2553 14843 2587
rect 14791 2515 14843 2553
rect 14911 2557 15016 2599
rect 14911 2523 14923 2557
rect 14957 2523 15016 2557
rect 14911 2515 15016 2523
rect 15046 2587 15096 2599
rect 15527 2599 15577 2643
rect 15255 2587 15373 2599
rect 15046 2563 15111 2587
rect 15046 2529 15056 2563
rect 15090 2529 15111 2563
rect 15046 2515 15111 2529
rect 15141 2563 15207 2587
rect 15141 2529 15163 2563
rect 15197 2529 15207 2563
rect 15141 2515 15207 2529
rect 15237 2515 15373 2587
rect 15403 2515 15445 2599
rect 15475 2561 15577 2599
rect 15475 2527 15509 2561
rect 15543 2527 15577 2561
rect 15475 2515 15577 2527
rect 15607 2587 15661 2643
rect 16257 2600 16309 2645
rect 15831 2587 15881 2599
rect 15607 2557 15676 2587
rect 15607 2523 15621 2557
rect 15655 2523 15676 2557
rect 15607 2515 15676 2523
rect 15706 2561 15785 2587
rect 15706 2527 15731 2561
rect 15765 2527 15785 2561
rect 15706 2515 15785 2527
rect 15815 2515 15881 2587
rect 15911 2557 16030 2599
rect 15911 2523 15943 2557
rect 15977 2523 16030 2557
rect 15911 2515 16030 2523
rect 16060 2515 16121 2599
rect 16151 2577 16203 2599
rect 16151 2543 16161 2577
rect 16195 2543 16203 2577
rect 16151 2515 16203 2543
rect 16257 2566 16265 2600
rect 16299 2566 16309 2600
rect 16257 2515 16309 2566
rect 16339 2633 16391 2645
rect 16339 2599 16349 2633
rect 16383 2599 16391 2633
rect 16542 2599 16594 2645
rect 16339 2565 16391 2599
rect 16339 2531 16349 2565
rect 16383 2531 16391 2565
rect 16339 2515 16391 2531
rect 16445 2587 16497 2599
rect 16445 2553 16453 2587
rect 16487 2553 16497 2587
rect 16445 2515 16497 2553
rect 16527 2581 16594 2599
rect 16527 2547 16550 2581
rect 16584 2547 16594 2581
rect 16527 2515 16594 2547
rect 16624 2611 16676 2645
rect 16624 2577 16634 2611
rect 16668 2577 16676 2611
rect 16624 2515 16676 2577
rect 17152 2322 17210 2334
rect 17152 2146 17164 2322
rect 17198 2146 17210 2322
rect 17152 2134 17210 2146
rect 17240 2322 17298 2334
rect 17240 2146 17252 2322
rect 17286 2146 17298 2322
rect 17240 2134 17298 2146
rect 160 1860 218 1872
rect 160 1684 172 1860
rect 206 1684 218 1860
rect 160 1672 218 1684
rect 418 1860 476 1872
rect 418 1684 430 1860
rect 464 1684 476 1860
rect 418 1672 476 1684
rect 540 1860 598 1872
rect 540 1684 552 1860
rect 586 1684 598 1860
rect 540 1672 598 1684
rect 798 1860 856 1872
rect 798 1684 810 1860
rect 844 1684 856 1860
rect 798 1672 856 1684
rect 920 1860 978 1872
rect 920 1684 932 1860
rect 966 1684 978 1860
rect 920 1672 978 1684
rect 1178 1860 1236 1872
rect 1178 1684 1190 1860
rect 1224 1684 1236 1860
rect 1178 1672 1236 1684
rect 1300 1860 1358 1872
rect 1300 1684 1312 1860
rect 1346 1684 1358 1860
rect 1300 1672 1358 1684
rect 1558 1860 1616 1872
rect 1558 1684 1570 1860
rect 1604 1684 1616 1860
rect 1558 1672 1616 1684
rect 1680 1860 1738 1872
rect 1680 1684 1692 1860
rect 1726 1684 1738 1860
rect 1680 1672 1738 1684
rect 1938 1860 1996 1872
rect 1938 1684 1950 1860
rect 1984 1684 1996 1860
rect 1938 1672 1996 1684
rect 2060 1860 2118 1872
rect 2060 1684 2072 1860
rect 2106 1684 2118 1860
rect 2060 1672 2118 1684
rect 2318 1860 2376 1872
rect 2318 1684 2330 1860
rect 2364 1684 2376 1860
rect 2318 1672 2376 1684
rect 2440 1860 2498 1872
rect 2440 1684 2452 1860
rect 2486 1684 2498 1860
rect 2440 1672 2498 1684
rect 2698 1860 2756 1872
rect 2698 1684 2710 1860
rect 2744 1684 2756 1860
rect 2698 1672 2756 1684
rect 2820 1860 2878 1872
rect 2820 1684 2832 1860
rect 2866 1684 2878 1860
rect 2820 1672 2878 1684
rect 3078 1860 3136 1872
rect 3078 1684 3090 1860
rect 3124 1684 3136 1860
rect 3078 1672 3136 1684
rect 160 1442 218 1454
rect 160 1266 172 1442
rect 206 1266 218 1442
rect 160 1254 218 1266
rect 418 1442 476 1454
rect 418 1266 430 1442
rect 464 1266 476 1442
rect 418 1254 476 1266
rect 540 1442 598 1454
rect 540 1266 552 1442
rect 586 1266 598 1442
rect 540 1254 598 1266
rect 798 1442 856 1454
rect 798 1266 810 1442
rect 844 1266 856 1442
rect 798 1254 856 1266
rect 920 1442 978 1454
rect 920 1266 932 1442
rect 966 1266 978 1442
rect 920 1254 978 1266
rect 1178 1442 1236 1454
rect 1178 1266 1190 1442
rect 1224 1266 1236 1442
rect 1178 1254 1236 1266
rect 1300 1442 1358 1454
rect 1300 1266 1312 1442
rect 1346 1266 1358 1442
rect 1300 1254 1358 1266
rect 1558 1442 1616 1454
rect 1558 1266 1570 1442
rect 1604 1266 1616 1442
rect 1558 1254 1616 1266
rect 1680 1442 1738 1454
rect 1680 1266 1692 1442
rect 1726 1266 1738 1442
rect 1680 1254 1738 1266
rect 1938 1442 1996 1454
rect 1938 1266 1950 1442
rect 1984 1266 1996 1442
rect 1938 1254 1996 1266
rect 2060 1442 2118 1454
rect 2060 1266 2072 1442
rect 2106 1266 2118 1442
rect 2060 1254 2118 1266
rect 2318 1442 2376 1454
rect 2318 1266 2330 1442
rect 2364 1266 2376 1442
rect 2318 1254 2376 1266
rect 2440 1442 2498 1454
rect 2440 1266 2452 1442
rect 2486 1266 2498 1442
rect 2440 1254 2498 1266
rect 2698 1442 2756 1454
rect 2698 1266 2710 1442
rect 2744 1266 2756 1442
rect 2698 1254 2756 1266
rect 2820 1442 2878 1454
rect 2820 1266 2832 1442
rect 2866 1266 2878 1442
rect 2820 1254 2878 1266
rect 3078 1442 3136 1454
rect 3078 1266 3090 1442
rect 3124 1266 3136 1442
rect 3078 1254 3136 1266
rect 160 1024 218 1036
rect 160 848 172 1024
rect 206 848 218 1024
rect 160 836 218 848
rect 418 1024 476 1036
rect 418 848 430 1024
rect 464 848 476 1024
rect 418 836 476 848
rect 540 1024 598 1036
rect 540 848 552 1024
rect 586 848 598 1024
rect 540 836 598 848
rect 798 1024 856 1036
rect 798 848 810 1024
rect 844 848 856 1024
rect 798 836 856 848
rect 920 1024 978 1036
rect 920 848 932 1024
rect 966 848 978 1024
rect 920 836 978 848
rect 1178 1024 1236 1036
rect 1178 848 1190 1024
rect 1224 848 1236 1024
rect 1178 836 1236 848
rect 1300 1024 1358 1036
rect 1300 848 1312 1024
rect 1346 848 1358 1024
rect 1300 836 1358 848
rect 1558 1024 1616 1036
rect 1558 848 1570 1024
rect 1604 848 1616 1024
rect 1558 836 1616 848
rect 1680 1024 1738 1036
rect 1680 848 1692 1024
rect 1726 848 1738 1024
rect 1680 836 1738 848
rect 1938 1024 1996 1036
rect 1938 848 1950 1024
rect 1984 848 1996 1024
rect 1938 836 1996 848
rect 2060 1024 2118 1036
rect 2060 848 2072 1024
rect 2106 848 2118 1024
rect 2060 836 2118 848
rect 2318 1024 2376 1036
rect 2318 848 2330 1024
rect 2364 848 2376 1024
rect 2318 836 2376 848
rect 2440 1024 2498 1036
rect 2440 848 2452 1024
rect 2486 848 2498 1024
rect 2440 836 2498 848
rect 2698 1024 2756 1036
rect 2698 848 2710 1024
rect 2744 848 2756 1024
rect 2698 836 2756 848
rect 2820 1024 2878 1036
rect 2820 848 2832 1024
rect 2866 848 2878 1024
rect 2820 836 2878 848
rect 3078 1024 3136 1036
rect 3078 848 3090 1024
rect 3124 848 3136 1024
rect 3078 836 3136 848
rect 160 606 218 618
rect 160 430 172 606
rect 206 430 218 606
rect 160 418 218 430
rect 418 606 476 618
rect 418 430 430 606
rect 464 430 476 606
rect 418 418 476 430
rect 540 606 598 618
rect 540 430 552 606
rect 586 430 598 606
rect 540 418 598 430
rect 798 606 856 618
rect 798 430 810 606
rect 844 430 856 606
rect 798 418 856 430
rect 920 606 978 618
rect 920 430 932 606
rect 966 430 978 606
rect 920 418 978 430
rect 1178 606 1236 618
rect 1178 430 1190 606
rect 1224 430 1236 606
rect 1178 418 1236 430
rect 1300 606 1358 618
rect 1300 430 1312 606
rect 1346 430 1358 606
rect 1300 418 1358 430
rect 1558 606 1616 618
rect 1558 430 1570 606
rect 1604 430 1616 606
rect 1558 418 1616 430
rect 1680 606 1738 618
rect 1680 430 1692 606
rect 1726 430 1738 606
rect 1680 418 1738 430
rect 1938 606 1996 618
rect 1938 430 1950 606
rect 1984 430 1996 606
rect 1938 418 1996 430
rect 2060 606 2118 618
rect 2060 430 2072 606
rect 2106 430 2118 606
rect 2060 418 2118 430
rect 2318 606 2376 618
rect 2318 430 2330 606
rect 2364 430 2376 606
rect 2318 418 2376 430
rect 2440 606 2498 618
rect 2440 430 2452 606
rect 2486 430 2498 606
rect 2440 418 2498 430
rect 2698 606 2756 618
rect 2698 430 2710 606
rect 2744 430 2756 606
rect 2698 418 2756 430
rect 2820 606 2878 618
rect 2820 430 2832 606
rect 2866 430 2878 606
rect 2820 418 2878 430
rect 3078 606 3136 618
rect 3078 430 3090 606
rect 3124 430 3136 606
rect 3078 418 3136 430
<< pdiff >>
rect 5796 5988 5854 6000
rect 5796 5812 5808 5988
rect 5842 5812 5854 5988
rect 5796 5800 5854 5812
rect 6054 5988 6112 6000
rect 6054 5812 6066 5988
rect 6100 5812 6112 5988
rect 6054 5800 6112 5812
rect 6312 5988 6370 6000
rect 6312 5812 6324 5988
rect 6358 5812 6370 5988
rect 6312 5800 6370 5812
rect 6570 5988 6628 6000
rect 6570 5812 6582 5988
rect 6616 5812 6628 5988
rect 6570 5800 6628 5812
rect 6828 5988 6886 6000
rect 6828 5812 6840 5988
rect 6874 5812 6886 5988
rect 6828 5800 6886 5812
rect 7086 5988 7144 6000
rect 7086 5812 7098 5988
rect 7132 5812 7144 5988
rect 7086 5800 7144 5812
rect 7344 5988 7402 6000
rect 7344 5812 7356 5988
rect 7390 5812 7402 5988
rect 7344 5800 7402 5812
rect 7456 5988 7514 6000
rect 7456 5812 7468 5988
rect 7502 5812 7514 5988
rect 7456 5800 7514 5812
rect 7714 5988 7772 6000
rect 7714 5812 7726 5988
rect 7760 5812 7772 5988
rect 7714 5800 7772 5812
rect 7836 5988 7894 6000
rect 7836 5812 7848 5988
rect 7882 5812 7894 5988
rect 7836 5800 7894 5812
rect 8094 5988 8152 6000
rect 8094 5812 8106 5988
rect 8140 5812 8152 5988
rect 8094 5800 8152 5812
rect 8352 5988 8410 6000
rect 8352 5812 8364 5988
rect 8398 5812 8410 5988
rect 8352 5800 8410 5812
rect 8610 5988 8668 6000
rect 8610 5812 8622 5988
rect 8656 5812 8668 5988
rect 8610 5800 8668 5812
rect 8868 5988 8926 6000
rect 8868 5812 8880 5988
rect 8914 5812 8926 5988
rect 8868 5800 8926 5812
rect 9126 5988 9184 6000
rect 9126 5812 9138 5988
rect 9172 5812 9184 5988
rect 9126 5800 9184 5812
rect 9256 5988 9314 6000
rect 9256 5812 9268 5988
rect 9302 5812 9314 5988
rect 9256 5800 9314 5812
rect 9514 5988 9572 6000
rect 9514 5812 9526 5988
rect 9560 5812 9572 5988
rect 9514 5800 9572 5812
rect 9772 5988 9830 6000
rect 9772 5812 9784 5988
rect 9818 5812 9830 5988
rect 9772 5800 9830 5812
rect 10030 5988 10088 6000
rect 10030 5812 10042 5988
rect 10076 5812 10088 5988
rect 10030 5800 10088 5812
rect 10288 5988 10346 6000
rect 10288 5812 10300 5988
rect 10334 5812 10346 5988
rect 10288 5800 10346 5812
rect 10546 5988 10604 6000
rect 10546 5812 10558 5988
rect 10592 5812 10604 5988
rect 10546 5800 10604 5812
rect 10676 5988 10734 6000
rect 10676 5812 10688 5988
rect 10722 5812 10734 5988
rect 10676 5800 10734 5812
rect 10934 5988 10992 6000
rect 10934 5812 10946 5988
rect 10980 5812 10992 5988
rect 10934 5800 10992 5812
rect 11056 5988 11114 6000
rect 11056 5812 11068 5988
rect 11102 5812 11114 5988
rect 11056 5800 11114 5812
rect 11314 5988 11372 6000
rect 11314 5812 11326 5988
rect 11360 5812 11372 5988
rect 11314 5800 11372 5812
rect 11572 5988 11630 6000
rect 11572 5812 11584 5988
rect 11618 5812 11630 5988
rect 11572 5800 11630 5812
rect 11830 5988 11888 6000
rect 11830 5812 11842 5988
rect 11876 5812 11888 5988
rect 11830 5800 11888 5812
rect 12088 5988 12146 6000
rect 12088 5812 12100 5988
rect 12134 5812 12146 5988
rect 12088 5800 12146 5812
rect 12346 5988 12404 6000
rect 12346 5812 12358 5988
rect 12392 5812 12404 5988
rect 12346 5800 12404 5812
rect 12604 5988 12662 6000
rect 12604 5812 12616 5988
rect 12650 5812 12662 5988
rect 12604 5800 12662 5812
rect 1756 4968 1814 4980
rect 1756 4592 1768 4968
rect 1802 4592 1814 4968
rect 1756 4580 1814 4592
rect 2014 4968 2072 4980
rect 2014 4592 2026 4968
rect 2060 4592 2072 4968
rect 2014 4580 2072 4592
rect 2136 4968 2194 4980
rect 2136 4592 2148 4968
rect 2182 4592 2194 4968
rect 2136 4580 2194 4592
rect 2394 4968 2452 4980
rect 2394 4592 2406 4968
rect 2440 4592 2452 4968
rect 2394 4580 2452 4592
rect 2516 4968 2574 4980
rect 2516 4592 2528 4968
rect 2562 4592 2574 4968
rect 2516 4580 2574 4592
rect 3574 4968 3632 4980
rect 3574 4592 3586 4968
rect 3620 4592 3632 4968
rect 3574 4580 3632 4592
rect 3696 4968 3754 4980
rect 3696 4592 3708 4968
rect 3742 4592 3754 4968
rect 3696 4580 3754 4592
rect 3954 4968 4012 4980
rect 3954 4592 3966 4968
rect 4000 4592 4012 4968
rect 3954 4580 4012 4592
rect 376 4288 434 4300
rect 376 3912 388 4288
rect 422 3912 434 4288
rect 376 3900 434 3912
rect 634 4288 692 4300
rect 634 3912 646 4288
rect 680 3912 692 4288
rect 634 3900 692 3912
rect 756 4288 814 4300
rect 756 3912 768 4288
rect 802 3912 814 4288
rect 756 3900 814 3912
rect 1014 4288 1072 4300
rect 1014 3912 1026 4288
rect 1060 3912 1072 4288
rect 1014 3900 1072 3912
rect 1272 4288 1330 4300
rect 1272 3912 1284 4288
rect 1318 3912 1330 4288
rect 1272 3900 1330 3912
rect 1396 4288 1454 4300
rect 1396 3912 1408 4288
rect 1442 3912 1454 4288
rect 1396 3900 1454 3912
rect 1654 4288 1712 4300
rect 1654 3912 1666 4288
rect 1700 3912 1712 4288
rect 1654 3900 1712 3912
rect 1912 4288 1970 4300
rect 1912 3912 1924 4288
rect 1958 3912 1970 4288
rect 1912 3900 1970 3912
rect 2170 4288 2228 4300
rect 2170 3912 2182 4288
rect 2216 3912 2228 4288
rect 2170 3900 2228 3912
rect 2428 4288 2486 4300
rect 2428 3912 2440 4288
rect 2474 3912 2486 4288
rect 2428 3900 2486 3912
rect 2556 4288 2614 4300
rect 2556 3912 2568 4288
rect 2602 3912 2614 4288
rect 2556 3900 2614 3912
rect 2814 4288 2872 4300
rect 2814 3912 2826 4288
rect 2860 3912 2872 4288
rect 2814 3900 2872 3912
rect 3072 4288 3130 4300
rect 3072 3912 3084 4288
rect 3118 3912 3130 4288
rect 3072 3900 3130 3912
rect 3330 4288 3388 4300
rect 3330 3912 3342 4288
rect 3376 3912 3388 4288
rect 3330 3900 3388 3912
rect 3588 4288 3646 4300
rect 3588 3912 3600 4288
rect 3634 3912 3646 4288
rect 3588 3900 3646 3912
rect 3716 4288 3774 4300
rect 3716 3912 3728 4288
rect 3762 3912 3774 4288
rect 3716 3900 3774 3912
rect 3974 4288 4032 4300
rect 3974 3912 3986 4288
rect 4020 3912 4032 4288
rect 3974 3900 4032 3912
rect 356 3048 414 3060
rect 356 2672 368 3048
rect 402 2672 414 3048
rect 356 2660 414 2672
rect 614 3048 672 3060
rect 614 2672 626 3048
rect 660 2672 672 3048
rect 614 2660 672 2672
rect 736 3048 794 3060
rect 736 2672 748 3048
rect 782 2672 794 3048
rect 736 2660 794 2672
rect 994 3048 1052 3060
rect 994 2672 1006 3048
rect 1040 2672 1052 3048
rect 994 2660 1052 2672
rect 1252 3048 1310 3060
rect 1252 2672 1264 3048
rect 1298 2672 1310 3048
rect 1252 2660 1310 2672
rect 1510 3048 1568 3060
rect 1510 2672 1522 3048
rect 1556 2672 1568 3048
rect 1510 2660 1568 2672
rect 1768 3048 1826 3060
rect 1768 2672 1780 3048
rect 1814 2672 1826 3048
rect 1768 2660 1826 2672
rect 2026 3048 2084 3060
rect 2026 2672 2038 3048
rect 2072 2672 2084 3048
rect 2026 2660 2084 2672
rect 2284 3048 2342 3060
rect 2284 2672 2296 3048
rect 2330 2672 2342 3048
rect 2284 2660 2342 2672
rect 2542 3048 2600 3060
rect 2542 2672 2554 3048
rect 2588 2672 2600 3048
rect 2542 2660 2600 2672
rect 2800 3048 2858 3060
rect 2800 2672 2812 3048
rect 2846 2672 2858 3048
rect 2800 2660 2858 2672
rect 2916 3048 2974 3060
rect 2916 2672 2928 3048
rect 2962 2672 2974 3048
rect 2916 2660 2974 2672
rect 3174 3048 3232 3060
rect 3174 2672 3186 3048
rect 3220 2672 3232 3048
rect 3174 2660 3232 2672
rect 14625 2945 14677 2959
rect 14625 2911 14633 2945
rect 14667 2911 14677 2945
rect 14625 2877 14677 2911
rect 14625 2843 14633 2877
rect 14667 2843 14677 2877
rect 14625 2831 14677 2843
rect 14707 2929 14761 2959
rect 14707 2895 14717 2929
rect 14751 2895 14761 2929
rect 14707 2831 14761 2895
rect 14791 2945 14843 2959
rect 14791 2911 14801 2945
rect 14835 2911 14843 2945
rect 14791 2877 14843 2911
rect 14976 2953 15028 2965
rect 14976 2919 14984 2953
rect 15018 2919 15028 2953
rect 14976 2881 15028 2919
rect 15058 2945 15120 2965
rect 15058 2911 15068 2945
rect 15102 2911 15120 2945
rect 15058 2881 15120 2911
rect 15150 2951 15219 2965
rect 15150 2917 15161 2951
rect 15195 2917 15219 2951
rect 15150 2881 15219 2917
rect 15249 2927 15359 2965
rect 15249 2893 15315 2927
rect 15349 2893 15359 2927
rect 15249 2881 15359 2893
rect 15389 2943 15456 2965
rect 15389 2909 15412 2943
rect 15446 2909 15456 2943
rect 15389 2881 15456 2909
rect 15486 2927 15538 2965
rect 15486 2893 15496 2927
rect 15530 2893 15538 2927
rect 15486 2881 15538 2893
rect 15601 2953 15653 2965
rect 15601 2919 15609 2953
rect 15643 2919 15653 2953
rect 14791 2843 14801 2877
rect 14835 2843 14843 2877
rect 14791 2831 14843 2843
rect 15601 2797 15653 2919
rect 15683 2945 15752 2965
rect 15683 2911 15697 2945
rect 15731 2911 15752 2945
rect 15683 2881 15752 2911
rect 15782 2952 15838 2965
rect 15782 2918 15794 2952
rect 15828 2918 15838 2952
rect 15782 2881 15838 2918
rect 15868 2881 15922 2965
rect 15952 2953 16030 2965
rect 15952 2919 15986 2953
rect 16020 2919 16030 2953
rect 15952 2881 16030 2919
rect 16060 2927 16114 2965
rect 16060 2893 16070 2927
rect 16104 2893 16114 2927
rect 16060 2881 16114 2893
rect 16144 2953 16278 2965
rect 16144 2919 16156 2953
rect 16190 2919 16234 2953
rect 16268 2919 16278 2953
rect 16144 2881 16278 2919
rect 15683 2797 15737 2881
rect 16228 2765 16278 2881
rect 16308 2945 16364 2965
rect 16308 2911 16318 2945
rect 16352 2911 16364 2945
rect 16308 2877 16364 2911
rect 16308 2843 16318 2877
rect 16352 2843 16364 2877
rect 16308 2809 16364 2843
rect 16445 2953 16497 2965
rect 16445 2919 16453 2953
rect 16487 2919 16497 2953
rect 16445 2885 16497 2919
rect 16445 2851 16453 2885
rect 16487 2851 16497 2885
rect 16445 2837 16497 2851
rect 16527 2953 16594 2965
rect 16527 2919 16550 2953
rect 16584 2919 16594 2953
rect 16527 2885 16594 2919
rect 16527 2851 16550 2885
rect 16584 2851 16594 2885
rect 16527 2837 16594 2851
rect 16308 2775 16318 2809
rect 16352 2775 16364 2809
rect 16308 2765 16364 2775
rect 16542 2817 16594 2837
rect 16542 2783 16550 2817
rect 16584 2783 16594 2817
rect 16542 2765 16594 2783
rect 16624 2917 16676 2965
rect 16624 2883 16634 2917
rect 16668 2883 16676 2917
rect 16624 2849 16676 2883
rect 16624 2815 16634 2849
rect 16668 2815 16676 2849
rect 16624 2765 16676 2815
rect 17152 3401 17210 3413
rect 17152 2825 17164 3401
rect 17198 2825 17210 3401
rect 17152 2813 17210 2825
rect 17240 3401 17298 3413
rect 17240 2825 17252 3401
rect 17286 2825 17298 3401
rect 17240 2813 17298 2825
<< ndiffc >>
rect 830 10562 864 10938
rect 918 10562 952 10938
rect 5838 4894 5872 5070
rect 6096 4894 6130 5070
rect 6354 4894 6388 5070
rect 6612 4894 6646 5070
rect 6870 4894 6904 5070
rect 7128 4894 7162 5070
rect 7386 4894 7420 5070
rect 7644 4894 7678 5070
rect 7902 4894 7936 5070
rect 8160 4894 8194 5070
rect 8418 4894 8452 5070
rect 8676 4894 8710 5070
rect 8934 4894 8968 5070
rect 9192 4894 9226 5070
rect 9450 4894 9484 5070
rect 9708 4894 9742 5070
rect 9966 4894 10000 5070
rect 10224 4894 10258 5070
rect 10482 4894 10516 5070
rect 10740 4894 10774 5070
rect 10998 4894 11032 5070
rect 11256 4894 11290 5070
rect 11514 4894 11548 5070
rect 5932 4060 5966 4236
rect 6190 4060 6224 4236
rect 6448 4060 6482 4236
rect 6706 4060 6740 4236
rect 6852 4060 6886 4236
rect 7110 4060 7144 4236
rect 7368 4060 7402 4236
rect 7626 4060 7660 4236
rect 7884 4060 7918 4236
rect 8142 4060 8176 4236
rect 8400 4060 8434 4236
rect 8658 4060 8692 4236
rect 8916 4060 8950 4236
rect 9174 4060 9208 4236
rect 9432 4060 9466 4236
rect 9690 4060 9724 4236
rect 9948 4060 9982 4236
rect 10206 4060 10240 4236
rect 10464 4060 10498 4236
rect 10722 4060 10756 4236
rect 10980 4060 11014 4236
rect 11238 4060 11272 4236
rect 11496 4060 11530 4236
rect 11754 4060 11788 4236
rect 12012 4060 12046 4236
rect 12270 4060 12304 4236
rect 14633 2553 14667 2587
rect 14717 2527 14751 2561
rect 14801 2553 14835 2587
rect 14923 2523 14957 2557
rect 15056 2529 15090 2563
rect 15163 2529 15197 2563
rect 15509 2527 15543 2561
rect 15621 2523 15655 2557
rect 15731 2527 15765 2561
rect 15943 2523 15977 2557
rect 16161 2543 16195 2577
rect 16265 2566 16299 2600
rect 16349 2599 16383 2633
rect 16349 2531 16383 2565
rect 16453 2553 16487 2587
rect 16550 2547 16584 2581
rect 16634 2577 16668 2611
rect 17164 2146 17198 2322
rect 17252 2146 17286 2322
rect 172 1684 206 1860
rect 430 1684 464 1860
rect 552 1684 586 1860
rect 810 1684 844 1860
rect 932 1684 966 1860
rect 1190 1684 1224 1860
rect 1312 1684 1346 1860
rect 1570 1684 1604 1860
rect 1692 1684 1726 1860
rect 1950 1684 1984 1860
rect 2072 1684 2106 1860
rect 2330 1684 2364 1860
rect 2452 1684 2486 1860
rect 2710 1684 2744 1860
rect 2832 1684 2866 1860
rect 3090 1684 3124 1860
rect 172 1266 206 1442
rect 430 1266 464 1442
rect 552 1266 586 1442
rect 810 1266 844 1442
rect 932 1266 966 1442
rect 1190 1266 1224 1442
rect 1312 1266 1346 1442
rect 1570 1266 1604 1442
rect 1692 1266 1726 1442
rect 1950 1266 1984 1442
rect 2072 1266 2106 1442
rect 2330 1266 2364 1442
rect 2452 1266 2486 1442
rect 2710 1266 2744 1442
rect 2832 1266 2866 1442
rect 3090 1266 3124 1442
rect 172 848 206 1024
rect 430 848 464 1024
rect 552 848 586 1024
rect 810 848 844 1024
rect 932 848 966 1024
rect 1190 848 1224 1024
rect 1312 848 1346 1024
rect 1570 848 1604 1024
rect 1692 848 1726 1024
rect 1950 848 1984 1024
rect 2072 848 2106 1024
rect 2330 848 2364 1024
rect 2452 848 2486 1024
rect 2710 848 2744 1024
rect 2832 848 2866 1024
rect 3090 848 3124 1024
rect 172 430 206 606
rect 430 430 464 606
rect 552 430 586 606
rect 810 430 844 606
rect 932 430 966 606
rect 1190 430 1224 606
rect 1312 430 1346 606
rect 1570 430 1604 606
rect 1692 430 1726 606
rect 1950 430 1984 606
rect 2072 430 2106 606
rect 2330 430 2364 606
rect 2452 430 2486 606
rect 2710 430 2744 606
rect 2832 430 2866 606
rect 3090 430 3124 606
<< pdiffc >>
rect 5808 5812 5842 5988
rect 6066 5812 6100 5988
rect 6324 5812 6358 5988
rect 6582 5812 6616 5988
rect 6840 5812 6874 5988
rect 7098 5812 7132 5988
rect 7356 5812 7390 5988
rect 7468 5812 7502 5988
rect 7726 5812 7760 5988
rect 7848 5812 7882 5988
rect 8106 5812 8140 5988
rect 8364 5812 8398 5988
rect 8622 5812 8656 5988
rect 8880 5812 8914 5988
rect 9138 5812 9172 5988
rect 9268 5812 9302 5988
rect 9526 5812 9560 5988
rect 9784 5812 9818 5988
rect 10042 5812 10076 5988
rect 10300 5812 10334 5988
rect 10558 5812 10592 5988
rect 10688 5812 10722 5988
rect 10946 5812 10980 5988
rect 11068 5812 11102 5988
rect 11326 5812 11360 5988
rect 11584 5812 11618 5988
rect 11842 5812 11876 5988
rect 12100 5812 12134 5988
rect 12358 5812 12392 5988
rect 12616 5812 12650 5988
rect 1768 4592 1802 4968
rect 2026 4592 2060 4968
rect 2148 4592 2182 4968
rect 2406 4592 2440 4968
rect 2528 4592 2562 4968
rect 3586 4592 3620 4968
rect 3708 4592 3742 4968
rect 3966 4592 4000 4968
rect 388 3912 422 4288
rect 646 3912 680 4288
rect 768 3912 802 4288
rect 1026 3912 1060 4288
rect 1284 3912 1318 4288
rect 1408 3912 1442 4288
rect 1666 3912 1700 4288
rect 1924 3912 1958 4288
rect 2182 3912 2216 4288
rect 2440 3912 2474 4288
rect 2568 3912 2602 4288
rect 2826 3912 2860 4288
rect 3084 3912 3118 4288
rect 3342 3912 3376 4288
rect 3600 3912 3634 4288
rect 3728 3912 3762 4288
rect 3986 3912 4020 4288
rect 368 2672 402 3048
rect 626 2672 660 3048
rect 748 2672 782 3048
rect 1006 2672 1040 3048
rect 1264 2672 1298 3048
rect 1522 2672 1556 3048
rect 1780 2672 1814 3048
rect 2038 2672 2072 3048
rect 2296 2672 2330 3048
rect 2554 2672 2588 3048
rect 2812 2672 2846 3048
rect 2928 2672 2962 3048
rect 3186 2672 3220 3048
rect 14633 2911 14667 2945
rect 14633 2843 14667 2877
rect 14717 2895 14751 2929
rect 14801 2911 14835 2945
rect 14984 2919 15018 2953
rect 15068 2911 15102 2945
rect 15161 2917 15195 2951
rect 15315 2893 15349 2927
rect 15412 2909 15446 2943
rect 15496 2893 15530 2927
rect 15609 2919 15643 2953
rect 14801 2843 14835 2877
rect 15697 2911 15731 2945
rect 15794 2918 15828 2952
rect 15986 2919 16020 2953
rect 16070 2893 16104 2927
rect 16156 2919 16190 2953
rect 16234 2919 16268 2953
rect 16318 2911 16352 2945
rect 16318 2843 16352 2877
rect 16453 2919 16487 2953
rect 16453 2851 16487 2885
rect 16550 2919 16584 2953
rect 16550 2851 16584 2885
rect 16318 2775 16352 2809
rect 16550 2783 16584 2817
rect 16634 2883 16668 2917
rect 16634 2815 16668 2849
rect 17164 2825 17198 3401
rect 17252 2825 17286 3401
<< psubdiff >>
rect 5996 31346 6092 31380
rect 6230 31346 6326 31380
rect 5996 31284 6030 31346
rect 6292 31284 6326 31346
rect 5996 29290 6030 29352
rect 6292 29290 6326 29352
rect 5996 29256 6092 29290
rect 6230 29256 6326 29290
rect 716 11090 812 11124
rect 970 11090 1066 11124
rect 716 11028 750 11090
rect 1032 11028 1066 11090
rect 716 10410 750 10472
rect 1032 10410 1066 10472
rect 716 10376 812 10410
rect 970 10376 1066 10410
rect 5736 5230 5832 5264
rect 11960 5230 12056 5264
rect 5736 5168 5770 5230
rect 12022 5168 12056 5230
rect 5736 4750 5770 4812
rect 12022 4750 12056 4812
rect 5736 4716 5832 4750
rect 11960 4716 12056 4750
rect 5816 4390 5912 4424
rect 12440 4390 12536 4424
rect 5816 4328 5850 4390
rect 12502 4328 12536 4390
rect 5816 3910 5850 3972
rect 12502 3910 12536 3972
rect 5816 3876 5912 3910
rect 12440 3876 12536 3910
rect 17050 2474 17146 2508
rect 17304 2474 17400 2508
rect 17050 2412 17084 2474
rect 17366 2412 17400 2474
rect 36 2010 132 2044
rect 3260 2010 3356 2044
rect 36 1948 70 2010
rect 3322 1948 3356 2010
rect 17050 1994 17084 2056
rect 17366 1994 17400 2056
rect 17050 1960 17146 1994
rect 17304 1960 17400 1994
rect 36 230 70 292
rect 3322 230 3356 292
rect 36 196 132 230
rect 3260 196 3356 230
<< nsubdiff >>
rect 5683 6183 5743 6217
rect 12717 6183 12777 6217
rect 5683 6157 5717 6183
rect 12743 6157 12777 6183
rect 5683 5637 5717 5663
rect 12743 5637 12777 5663
rect 5683 5603 5743 5637
rect 12717 5603 12777 5637
rect 243 5223 303 5257
rect 4137 5223 4197 5257
rect 243 5197 277 5223
rect 4163 5197 4197 5223
rect 243 3697 277 3723
rect 4163 3697 4197 3723
rect 243 3663 303 3697
rect 4137 3663 4197 3697
rect 17050 3562 17146 3596
rect 17304 3562 17400 3596
rect 17050 3500 17084 3562
rect 203 3303 263 3337
rect 3297 3303 3357 3337
rect 203 3277 237 3303
rect 3323 3277 3357 3303
rect 203 2377 237 2403
rect 14420 2950 14520 2970
rect 14420 2910 14450 2950
rect 14490 2910 14520 2950
rect 14420 2880 14520 2910
rect 17366 3500 17400 3562
rect 17050 2664 17084 2726
rect 17366 2664 17400 2726
rect 17050 2630 17146 2664
rect 17304 2630 17400 2664
rect 3323 2377 3357 2403
rect 203 2343 263 2377
rect 3297 2343 3357 2377
<< psubdiffcont >>
rect 6092 31346 6230 31380
rect 5996 29352 6030 31284
rect 6292 29352 6326 31284
rect 6092 29256 6230 29290
rect 812 11090 970 11124
rect 716 10472 750 11028
rect 1032 10472 1066 11028
rect 812 10376 970 10410
rect 5832 5230 11960 5264
rect 5736 4812 5770 5168
rect 12022 4812 12056 5168
rect 5832 4716 11960 4750
rect 5912 4390 12440 4424
rect 5816 3972 5850 4328
rect 12502 3972 12536 4328
rect 5912 3876 12440 3910
rect 17146 2474 17304 2508
rect 17050 2056 17084 2412
rect 132 2010 3260 2044
rect 36 292 70 1948
rect 17366 2056 17400 2412
rect 17146 1960 17304 1994
rect 3322 292 3356 1948
rect 132 196 3260 230
<< nsubdiffcont >>
rect 5743 6183 12717 6217
rect 5683 5663 5717 6157
rect 12743 5663 12777 6157
rect 5743 5603 12717 5637
rect 303 5223 4137 5257
rect 243 3723 277 5197
rect 4163 3723 4197 5197
rect 303 3663 4137 3697
rect 17146 3562 17304 3596
rect 263 3303 3297 3337
rect 203 2403 237 3277
rect 3323 2403 3357 3277
rect 14450 2910 14490 2950
rect 17050 2726 17084 3500
rect 17366 2726 17400 3500
rect 17146 2630 17304 2664
rect 263 2343 3297 2377
<< poly >>
rect 858 11022 924 11038
rect 858 10988 874 11022
rect 908 10988 924 11022
rect 858 10972 924 10988
rect 876 10950 906 10972
rect 876 10528 906 10550
rect 858 10512 924 10528
rect 858 10478 874 10512
rect 908 10478 924 10512
rect 858 10462 924 10478
rect 5854 6081 6054 6097
rect 5854 6047 5870 6081
rect 6038 6047 6054 6081
rect 5854 6000 6054 6047
rect 6112 6081 6312 6097
rect 6112 6047 6128 6081
rect 6296 6047 6312 6081
rect 6112 6000 6312 6047
rect 6370 6081 6570 6097
rect 6370 6047 6386 6081
rect 6554 6047 6570 6081
rect 6370 6000 6570 6047
rect 6628 6081 6828 6097
rect 6628 6047 6644 6081
rect 6812 6047 6828 6081
rect 6628 6000 6828 6047
rect 6886 6081 7086 6097
rect 6886 6047 6902 6081
rect 7070 6047 7086 6081
rect 6886 6000 7086 6047
rect 7144 6081 7344 6097
rect 7144 6047 7160 6081
rect 7328 6047 7344 6081
rect 7144 6000 7344 6047
rect 7514 6081 7714 6097
rect 7514 6047 7530 6081
rect 7698 6047 7714 6081
rect 7514 6000 7714 6047
rect 7894 6081 8094 6097
rect 7894 6047 7910 6081
rect 8078 6047 8094 6081
rect 7894 6000 8094 6047
rect 8152 6081 8352 6097
rect 8152 6047 8168 6081
rect 8336 6047 8352 6081
rect 8152 6000 8352 6047
rect 8410 6081 8610 6097
rect 8410 6047 8426 6081
rect 8594 6047 8610 6081
rect 8410 6000 8610 6047
rect 8668 6081 8868 6097
rect 8668 6047 8684 6081
rect 8852 6047 8868 6081
rect 8668 6000 8868 6047
rect 8926 6081 9126 6097
rect 8926 6047 8942 6081
rect 9110 6047 9126 6081
rect 8926 6000 9126 6047
rect 9314 6081 9514 6097
rect 9314 6047 9330 6081
rect 9498 6047 9514 6081
rect 9314 6000 9514 6047
rect 9572 6081 9772 6097
rect 9572 6047 9588 6081
rect 9756 6047 9772 6081
rect 9572 6000 9772 6047
rect 9830 6081 10030 6097
rect 9830 6047 9846 6081
rect 10014 6047 10030 6081
rect 9830 6000 10030 6047
rect 10088 6081 10288 6097
rect 10088 6047 10104 6081
rect 10272 6047 10288 6081
rect 10088 6000 10288 6047
rect 10346 6081 10546 6097
rect 10346 6047 10362 6081
rect 10530 6047 10546 6081
rect 10346 6000 10546 6047
rect 10734 6081 10934 6097
rect 10734 6047 10750 6081
rect 10918 6047 10934 6081
rect 10734 6000 10934 6047
rect 11114 6081 11314 6097
rect 11114 6047 11130 6081
rect 11298 6047 11314 6081
rect 11114 6000 11314 6047
rect 11372 6081 11572 6097
rect 11372 6047 11388 6081
rect 11556 6047 11572 6081
rect 11372 6000 11572 6047
rect 11630 6081 11830 6097
rect 11630 6047 11646 6081
rect 11814 6047 11830 6081
rect 11630 6000 11830 6047
rect 11888 6081 12088 6097
rect 11888 6047 11904 6081
rect 12072 6047 12088 6081
rect 11888 6000 12088 6047
rect 12146 6081 12346 6097
rect 12146 6047 12162 6081
rect 12330 6047 12346 6081
rect 12146 6000 12346 6047
rect 12404 6081 12604 6097
rect 12404 6047 12420 6081
rect 12588 6047 12604 6081
rect 12404 6000 12604 6047
rect 5854 5753 6054 5800
rect 5854 5719 5870 5753
rect 6038 5719 6054 5753
rect 5854 5703 6054 5719
rect 6112 5753 6312 5800
rect 6112 5719 6128 5753
rect 6296 5719 6312 5753
rect 6112 5703 6312 5719
rect 6370 5753 6570 5800
rect 6370 5719 6386 5753
rect 6554 5719 6570 5753
rect 6370 5703 6570 5719
rect 6628 5753 6828 5800
rect 6628 5719 6644 5753
rect 6812 5719 6828 5753
rect 6628 5703 6828 5719
rect 6886 5753 7086 5800
rect 6886 5719 6902 5753
rect 7070 5719 7086 5753
rect 6886 5703 7086 5719
rect 7144 5753 7344 5800
rect 7144 5719 7160 5753
rect 7328 5719 7344 5753
rect 7144 5703 7344 5719
rect 7514 5753 7714 5800
rect 7514 5719 7530 5753
rect 7698 5719 7714 5753
rect 7514 5703 7714 5719
rect 7894 5753 8094 5800
rect 7894 5719 7910 5753
rect 8078 5719 8094 5753
rect 7894 5703 8094 5719
rect 8152 5753 8352 5800
rect 8152 5719 8168 5753
rect 8336 5719 8352 5753
rect 8152 5703 8352 5719
rect 8410 5753 8610 5800
rect 8410 5719 8426 5753
rect 8594 5719 8610 5753
rect 8410 5703 8610 5719
rect 8668 5753 8868 5800
rect 8668 5719 8684 5753
rect 8852 5719 8868 5753
rect 8668 5703 8868 5719
rect 8926 5753 9126 5800
rect 8926 5719 8942 5753
rect 9110 5719 9126 5753
rect 8926 5703 9126 5719
rect 9314 5753 9514 5800
rect 9314 5719 9330 5753
rect 9498 5719 9514 5753
rect 9314 5703 9514 5719
rect 9572 5753 9772 5800
rect 9572 5719 9588 5753
rect 9756 5719 9772 5753
rect 9572 5703 9772 5719
rect 9830 5753 10030 5800
rect 9830 5719 9846 5753
rect 10014 5719 10030 5753
rect 9830 5703 10030 5719
rect 10088 5753 10288 5800
rect 10088 5719 10104 5753
rect 10272 5719 10288 5753
rect 10088 5703 10288 5719
rect 10346 5753 10546 5800
rect 10346 5719 10362 5753
rect 10530 5719 10546 5753
rect 10346 5703 10546 5719
rect 10734 5753 10934 5800
rect 10734 5719 10750 5753
rect 10918 5719 10934 5753
rect 10734 5703 10934 5719
rect 11114 5753 11314 5800
rect 11114 5719 11130 5753
rect 11298 5719 11314 5753
rect 11114 5703 11314 5719
rect 11372 5753 11572 5800
rect 11372 5719 11388 5753
rect 11556 5719 11572 5753
rect 11372 5703 11572 5719
rect 11630 5753 11830 5800
rect 11630 5719 11646 5753
rect 11814 5719 11830 5753
rect 11630 5703 11830 5719
rect 11888 5753 12088 5800
rect 11888 5719 11904 5753
rect 12072 5719 12088 5753
rect 11888 5703 12088 5719
rect 12146 5753 12346 5800
rect 12146 5719 12162 5753
rect 12330 5719 12346 5753
rect 12146 5703 12346 5719
rect 12404 5753 12604 5800
rect 12404 5719 12420 5753
rect 12588 5719 12604 5753
rect 12404 5703 12604 5719
rect 1814 5061 2014 5077
rect 1814 5027 1830 5061
rect 1998 5027 2014 5061
rect 1814 4980 2014 5027
rect 2194 5061 2394 5077
rect 2194 5027 2210 5061
rect 2378 5027 2394 5061
rect 2194 4980 2394 5027
rect 2574 5061 3574 5077
rect 2574 5027 2590 5061
rect 3558 5027 3574 5061
rect 2574 4980 3574 5027
rect 3754 5061 3954 5077
rect 3754 5027 3770 5061
rect 3938 5027 3954 5061
rect 3754 4980 3954 5027
rect 1814 4533 2014 4580
rect 1814 4499 1830 4533
rect 1998 4499 2014 4533
rect 1814 4483 2014 4499
rect 2194 4533 2394 4580
rect 2194 4499 2210 4533
rect 2378 4499 2394 4533
rect 2194 4483 2394 4499
rect 2574 4533 3574 4580
rect 2574 4499 2590 4533
rect 3558 4499 3574 4533
rect 2574 4483 3574 4499
rect 3754 4533 3954 4580
rect 3754 4499 3770 4533
rect 3938 4499 3954 4533
rect 3754 4483 3954 4499
rect 434 4381 634 4397
rect 434 4347 450 4381
rect 618 4347 634 4381
rect 434 4300 634 4347
rect 814 4381 1014 4397
rect 814 4347 830 4381
rect 998 4347 1014 4381
rect 814 4300 1014 4347
rect 1072 4381 1272 4397
rect 1072 4347 1088 4381
rect 1256 4347 1272 4381
rect 1072 4300 1272 4347
rect 1454 4381 1654 4397
rect 1454 4347 1470 4381
rect 1638 4347 1654 4381
rect 1454 4300 1654 4347
rect 1712 4381 1912 4397
rect 1712 4347 1728 4381
rect 1896 4347 1912 4381
rect 1712 4300 1912 4347
rect 1970 4381 2170 4397
rect 1970 4347 1986 4381
rect 2154 4347 2170 4381
rect 1970 4300 2170 4347
rect 2228 4381 2428 4397
rect 2228 4347 2244 4381
rect 2412 4347 2428 4381
rect 2228 4300 2428 4347
rect 2614 4381 2814 4397
rect 2614 4347 2630 4381
rect 2798 4347 2814 4381
rect 2614 4300 2814 4347
rect 2872 4381 3072 4397
rect 2872 4347 2888 4381
rect 3056 4347 3072 4381
rect 2872 4300 3072 4347
rect 3130 4381 3330 4397
rect 3130 4347 3146 4381
rect 3314 4347 3330 4381
rect 3130 4300 3330 4347
rect 3388 4381 3588 4397
rect 3388 4347 3404 4381
rect 3572 4347 3588 4381
rect 3388 4300 3588 4347
rect 3774 4381 3974 4397
rect 3774 4347 3790 4381
rect 3958 4347 3974 4381
rect 3774 4300 3974 4347
rect 434 3853 634 3900
rect 434 3819 450 3853
rect 618 3819 634 3853
rect 434 3803 634 3819
rect 814 3853 1014 3900
rect 814 3819 830 3853
rect 998 3819 1014 3853
rect 814 3803 1014 3819
rect 1072 3853 1272 3900
rect 1072 3819 1088 3853
rect 1256 3819 1272 3853
rect 1072 3803 1272 3819
rect 1454 3853 1654 3900
rect 1454 3819 1470 3853
rect 1638 3819 1654 3853
rect 1454 3803 1654 3819
rect 1712 3853 1912 3900
rect 1712 3819 1728 3853
rect 1896 3819 1912 3853
rect 1712 3803 1912 3819
rect 1970 3853 2170 3900
rect 1970 3819 1986 3853
rect 2154 3819 2170 3853
rect 1970 3803 2170 3819
rect 2228 3853 2428 3900
rect 2228 3819 2244 3853
rect 2412 3819 2428 3853
rect 2228 3803 2428 3819
rect 2614 3853 2814 3900
rect 2614 3819 2630 3853
rect 2798 3819 2814 3853
rect 2614 3803 2814 3819
rect 2872 3853 3072 3900
rect 2872 3819 2888 3853
rect 3056 3819 3072 3853
rect 2872 3803 3072 3819
rect 3130 3853 3330 3900
rect 3130 3819 3146 3853
rect 3314 3819 3330 3853
rect 3130 3803 3330 3819
rect 3388 3853 3588 3900
rect 3388 3819 3404 3853
rect 3572 3819 3588 3853
rect 3388 3803 3588 3819
rect 3774 3853 3974 3900
rect 3774 3819 3790 3853
rect 3958 3819 3974 3853
rect 3774 3803 3974 3819
rect 5884 5154 6084 5170
rect 5884 5120 5900 5154
rect 6068 5120 6084 5154
rect 5884 5082 6084 5120
rect 6142 5154 6342 5170
rect 6142 5120 6158 5154
rect 6326 5120 6342 5154
rect 6142 5082 6342 5120
rect 6400 5154 6600 5170
rect 6400 5120 6416 5154
rect 6584 5120 6600 5154
rect 6400 5082 6600 5120
rect 6658 5154 6858 5170
rect 6658 5120 6674 5154
rect 6842 5120 6858 5154
rect 6658 5082 6858 5120
rect 6916 5154 7116 5170
rect 6916 5120 6932 5154
rect 7100 5120 7116 5154
rect 6916 5082 7116 5120
rect 7174 5154 7374 5170
rect 7174 5120 7190 5154
rect 7358 5120 7374 5154
rect 7174 5082 7374 5120
rect 7432 5154 7632 5170
rect 7432 5120 7448 5154
rect 7616 5120 7632 5154
rect 7432 5082 7632 5120
rect 7690 5154 7890 5170
rect 7690 5120 7706 5154
rect 7874 5120 7890 5154
rect 7690 5082 7890 5120
rect 7948 5154 8148 5170
rect 7948 5120 7964 5154
rect 8132 5120 8148 5154
rect 7948 5082 8148 5120
rect 8206 5154 8406 5170
rect 8206 5120 8222 5154
rect 8390 5120 8406 5154
rect 8206 5082 8406 5120
rect 8464 5154 8664 5170
rect 8464 5120 8480 5154
rect 8648 5120 8664 5154
rect 8464 5082 8664 5120
rect 8722 5154 8922 5170
rect 8722 5120 8738 5154
rect 8906 5120 8922 5154
rect 8722 5082 8922 5120
rect 8980 5154 9180 5170
rect 8980 5120 8996 5154
rect 9164 5120 9180 5154
rect 8980 5082 9180 5120
rect 9238 5154 9438 5170
rect 9238 5120 9254 5154
rect 9422 5120 9438 5154
rect 9238 5082 9438 5120
rect 9496 5154 9696 5170
rect 9496 5120 9512 5154
rect 9680 5120 9696 5154
rect 9496 5082 9696 5120
rect 9754 5154 9954 5170
rect 9754 5120 9770 5154
rect 9938 5120 9954 5154
rect 9754 5082 9954 5120
rect 10012 5154 10212 5170
rect 10012 5120 10028 5154
rect 10196 5120 10212 5154
rect 10012 5082 10212 5120
rect 10270 5154 10470 5170
rect 10270 5120 10286 5154
rect 10454 5120 10470 5154
rect 10270 5082 10470 5120
rect 10528 5154 10728 5170
rect 10528 5120 10544 5154
rect 10712 5120 10728 5154
rect 10528 5082 10728 5120
rect 10786 5154 10986 5170
rect 10786 5120 10802 5154
rect 10970 5120 10986 5154
rect 10786 5082 10986 5120
rect 11044 5154 11244 5170
rect 11044 5120 11060 5154
rect 11228 5120 11244 5154
rect 11044 5082 11244 5120
rect 11302 5154 11502 5170
rect 11302 5120 11318 5154
rect 11486 5120 11502 5154
rect 11302 5082 11502 5120
rect 5884 4844 6084 4882
rect 5884 4810 5900 4844
rect 6068 4810 6084 4844
rect 5884 4794 6084 4810
rect 6142 4844 6342 4882
rect 6142 4810 6158 4844
rect 6326 4810 6342 4844
rect 6142 4794 6342 4810
rect 6400 4844 6600 4882
rect 6400 4810 6416 4844
rect 6584 4810 6600 4844
rect 6400 4794 6600 4810
rect 6658 4844 6858 4882
rect 6658 4810 6674 4844
rect 6842 4810 6858 4844
rect 6658 4794 6858 4810
rect 6916 4844 7116 4882
rect 6916 4810 6932 4844
rect 7100 4810 7116 4844
rect 6916 4794 7116 4810
rect 7174 4844 7374 4882
rect 7174 4810 7190 4844
rect 7358 4810 7374 4844
rect 7174 4794 7374 4810
rect 7432 4844 7632 4882
rect 7432 4810 7448 4844
rect 7616 4810 7632 4844
rect 7432 4794 7632 4810
rect 7690 4844 7890 4882
rect 7690 4810 7706 4844
rect 7874 4810 7890 4844
rect 7690 4794 7890 4810
rect 7948 4844 8148 4882
rect 7948 4810 7964 4844
rect 8132 4810 8148 4844
rect 7948 4794 8148 4810
rect 8206 4844 8406 4882
rect 8206 4810 8222 4844
rect 8390 4810 8406 4844
rect 8206 4794 8406 4810
rect 8464 4844 8664 4882
rect 8464 4810 8480 4844
rect 8648 4810 8664 4844
rect 8464 4794 8664 4810
rect 8722 4844 8922 4882
rect 8722 4810 8738 4844
rect 8906 4810 8922 4844
rect 8722 4794 8922 4810
rect 8980 4844 9180 4882
rect 8980 4810 8996 4844
rect 9164 4810 9180 4844
rect 8980 4794 9180 4810
rect 9238 4844 9438 4882
rect 9238 4810 9254 4844
rect 9422 4810 9438 4844
rect 9238 4794 9438 4810
rect 9496 4844 9696 4882
rect 9496 4810 9512 4844
rect 9680 4810 9696 4844
rect 9496 4794 9696 4810
rect 9754 4844 9954 4882
rect 9754 4810 9770 4844
rect 9938 4810 9954 4844
rect 9754 4794 9954 4810
rect 10012 4844 10212 4882
rect 10012 4810 10028 4844
rect 10196 4810 10212 4844
rect 10012 4794 10212 4810
rect 10270 4844 10470 4882
rect 10270 4810 10286 4844
rect 10454 4810 10470 4844
rect 10270 4794 10470 4810
rect 10528 4844 10728 4882
rect 10528 4810 10544 4844
rect 10712 4810 10728 4844
rect 10528 4794 10728 4810
rect 10786 4844 10986 4882
rect 10786 4810 10802 4844
rect 10970 4810 10986 4844
rect 10786 4794 10986 4810
rect 11044 4844 11244 4882
rect 11044 4810 11060 4844
rect 11228 4810 11244 4844
rect 11044 4794 11244 4810
rect 11302 4844 11502 4882
rect 11302 4810 11318 4844
rect 11486 4810 11502 4844
rect 11302 4794 11502 4810
rect 5978 4320 6178 4336
rect 5978 4286 5994 4320
rect 6162 4286 6178 4320
rect 5978 4248 6178 4286
rect 6236 4320 6436 4336
rect 6236 4286 6252 4320
rect 6420 4286 6436 4320
rect 6236 4248 6436 4286
rect 6494 4320 6694 4336
rect 6494 4286 6510 4320
rect 6678 4286 6694 4320
rect 6494 4248 6694 4286
rect 6898 4320 7098 4336
rect 6898 4286 6914 4320
rect 7082 4286 7098 4320
rect 6898 4248 7098 4286
rect 7156 4320 7356 4336
rect 7156 4286 7172 4320
rect 7340 4286 7356 4320
rect 7156 4248 7356 4286
rect 7414 4320 7614 4336
rect 7414 4286 7430 4320
rect 7598 4286 7614 4320
rect 7414 4248 7614 4286
rect 7672 4320 7872 4336
rect 7672 4286 7688 4320
rect 7856 4286 7872 4320
rect 7672 4248 7872 4286
rect 7930 4320 8130 4336
rect 7930 4286 7946 4320
rect 8114 4286 8130 4320
rect 7930 4248 8130 4286
rect 8188 4320 8388 4336
rect 8188 4286 8204 4320
rect 8372 4286 8388 4320
rect 8188 4248 8388 4286
rect 8446 4320 8646 4336
rect 8446 4286 8462 4320
rect 8630 4286 8646 4320
rect 8446 4248 8646 4286
rect 8704 4320 8904 4336
rect 8704 4286 8720 4320
rect 8888 4286 8904 4320
rect 8704 4248 8904 4286
rect 8962 4320 9162 4336
rect 8962 4286 8978 4320
rect 9146 4286 9162 4320
rect 8962 4248 9162 4286
rect 9220 4320 9420 4336
rect 9220 4286 9236 4320
rect 9404 4286 9420 4320
rect 9220 4248 9420 4286
rect 9478 4320 9678 4336
rect 9478 4286 9494 4320
rect 9662 4286 9678 4320
rect 9478 4248 9678 4286
rect 9736 4320 9936 4336
rect 9736 4286 9752 4320
rect 9920 4286 9936 4320
rect 9736 4248 9936 4286
rect 9994 4320 10194 4336
rect 9994 4286 10010 4320
rect 10178 4286 10194 4320
rect 9994 4248 10194 4286
rect 10252 4320 10452 4336
rect 10252 4286 10268 4320
rect 10436 4286 10452 4320
rect 10252 4248 10452 4286
rect 10510 4320 10710 4336
rect 10510 4286 10526 4320
rect 10694 4286 10710 4320
rect 10510 4248 10710 4286
rect 10768 4320 10968 4336
rect 10768 4286 10784 4320
rect 10952 4286 10968 4320
rect 10768 4248 10968 4286
rect 11026 4320 11226 4336
rect 11026 4286 11042 4320
rect 11210 4286 11226 4320
rect 11026 4248 11226 4286
rect 11284 4320 11484 4336
rect 11284 4286 11300 4320
rect 11468 4286 11484 4320
rect 11284 4248 11484 4286
rect 11542 4320 11742 4336
rect 11542 4286 11558 4320
rect 11726 4286 11742 4320
rect 11542 4248 11742 4286
rect 11800 4320 12000 4336
rect 11800 4286 11816 4320
rect 11984 4286 12000 4320
rect 11800 4248 12000 4286
rect 12058 4320 12258 4336
rect 12058 4286 12074 4320
rect 12242 4286 12258 4320
rect 12058 4248 12258 4286
rect 5978 4010 6178 4048
rect 5978 3976 5994 4010
rect 6162 3976 6178 4010
rect 5978 3960 6178 3976
rect 6236 4010 6436 4048
rect 6236 3976 6252 4010
rect 6420 3976 6436 4010
rect 6236 3960 6436 3976
rect 6494 4010 6694 4048
rect 6494 3976 6510 4010
rect 6678 3976 6694 4010
rect 6494 3960 6694 3976
rect 6898 4010 7098 4048
rect 6898 3976 6914 4010
rect 7082 3976 7098 4010
rect 6898 3960 7098 3976
rect 7156 4010 7356 4048
rect 7156 3976 7172 4010
rect 7340 3976 7356 4010
rect 7156 3960 7356 3976
rect 7414 4010 7614 4048
rect 7414 3976 7430 4010
rect 7598 3976 7614 4010
rect 7414 3960 7614 3976
rect 7672 4010 7872 4048
rect 7672 3976 7688 4010
rect 7856 3976 7872 4010
rect 7672 3960 7872 3976
rect 7930 4010 8130 4048
rect 7930 3976 7946 4010
rect 8114 3976 8130 4010
rect 7930 3960 8130 3976
rect 8188 4010 8388 4048
rect 8188 3976 8204 4010
rect 8372 3976 8388 4010
rect 8188 3960 8388 3976
rect 8446 4010 8646 4048
rect 8446 3976 8462 4010
rect 8630 3976 8646 4010
rect 8446 3960 8646 3976
rect 8704 4010 8904 4048
rect 8704 3976 8720 4010
rect 8888 3976 8904 4010
rect 8704 3960 8904 3976
rect 8962 4010 9162 4048
rect 8962 3976 8978 4010
rect 9146 3976 9162 4010
rect 8962 3960 9162 3976
rect 9220 4010 9420 4048
rect 9220 3976 9236 4010
rect 9404 3976 9420 4010
rect 9220 3960 9420 3976
rect 9478 4010 9678 4048
rect 9478 3976 9494 4010
rect 9662 3976 9678 4010
rect 9478 3960 9678 3976
rect 9736 4010 9936 4048
rect 9736 3976 9752 4010
rect 9920 3976 9936 4010
rect 9736 3960 9936 3976
rect 9994 4010 10194 4048
rect 9994 3976 10010 4010
rect 10178 3976 10194 4010
rect 9994 3960 10194 3976
rect 10252 4010 10452 4048
rect 10252 3976 10268 4010
rect 10436 3976 10452 4010
rect 10252 3960 10452 3976
rect 10510 4010 10710 4048
rect 10510 3976 10526 4010
rect 10694 3976 10710 4010
rect 10510 3960 10710 3976
rect 10768 4010 10968 4048
rect 10768 3976 10784 4010
rect 10952 3976 10968 4010
rect 10768 3960 10968 3976
rect 11026 4010 11226 4048
rect 11026 3976 11042 4010
rect 11210 3976 11226 4010
rect 11026 3960 11226 3976
rect 11284 4010 11484 4048
rect 11284 3976 11300 4010
rect 11468 3976 11484 4010
rect 11284 3960 11484 3976
rect 11542 4010 11742 4048
rect 11542 3976 11558 4010
rect 11726 3976 11742 4010
rect 11542 3960 11742 3976
rect 11800 4010 12000 4048
rect 11800 3976 11816 4010
rect 11984 3976 12000 4010
rect 11800 3960 12000 3976
rect 12058 4010 12258 4048
rect 12058 3976 12074 4010
rect 12242 3976 12258 4010
rect 12058 3960 12258 3976
rect 414 3141 614 3157
rect 414 3107 430 3141
rect 598 3107 614 3141
rect 414 3060 614 3107
rect 794 3141 994 3157
rect 794 3107 810 3141
rect 978 3107 994 3141
rect 794 3060 994 3107
rect 1052 3141 1252 3157
rect 1052 3107 1068 3141
rect 1236 3107 1252 3141
rect 1052 3060 1252 3107
rect 1310 3141 1510 3157
rect 1310 3107 1326 3141
rect 1494 3107 1510 3141
rect 1310 3060 1510 3107
rect 1568 3141 1768 3157
rect 1568 3107 1584 3141
rect 1752 3107 1768 3141
rect 1568 3060 1768 3107
rect 1826 3141 2026 3157
rect 1826 3107 1842 3141
rect 2010 3107 2026 3141
rect 1826 3060 2026 3107
rect 2084 3141 2284 3157
rect 2084 3107 2100 3141
rect 2268 3107 2284 3141
rect 2084 3060 2284 3107
rect 2342 3141 2542 3157
rect 2342 3107 2358 3141
rect 2526 3107 2542 3141
rect 2342 3060 2542 3107
rect 2600 3141 2800 3157
rect 2600 3107 2616 3141
rect 2784 3107 2800 3141
rect 2600 3060 2800 3107
rect 2974 3141 3174 3157
rect 2974 3107 2990 3141
rect 3158 3107 3174 3141
rect 2974 3060 3174 3107
rect 414 2613 614 2660
rect 414 2579 430 2613
rect 598 2579 614 2613
rect 414 2563 614 2579
rect 794 2613 994 2660
rect 794 2579 810 2613
rect 978 2579 994 2613
rect 794 2563 994 2579
rect 1052 2613 1252 2660
rect 1052 2579 1068 2613
rect 1236 2579 1252 2613
rect 1052 2563 1252 2579
rect 1310 2613 1510 2660
rect 1310 2579 1326 2613
rect 1494 2579 1510 2613
rect 1310 2563 1510 2579
rect 1568 2613 1768 2660
rect 1568 2579 1584 2613
rect 1752 2579 1768 2613
rect 1568 2563 1768 2579
rect 1826 2613 2026 2660
rect 1826 2579 1842 2613
rect 2010 2579 2026 2613
rect 1826 2563 2026 2579
rect 2084 2613 2284 2660
rect 2084 2579 2100 2613
rect 2268 2579 2284 2613
rect 2084 2563 2284 2579
rect 2342 2613 2542 2660
rect 2342 2579 2358 2613
rect 2526 2579 2542 2613
rect 2342 2563 2542 2579
rect 2600 2613 2800 2660
rect 2600 2579 2616 2613
rect 2784 2579 2800 2613
rect 2600 2563 2800 2579
rect 2974 2613 3174 2660
rect 2974 2579 2990 2613
rect 3158 2579 3174 2613
rect 2974 2563 3174 2579
rect 14677 2959 14707 2985
rect 14761 2959 14791 2985
rect 15028 2965 15058 2991
rect 15120 2965 15150 2991
rect 15219 2965 15249 2991
rect 15359 2965 15389 2991
rect 15456 2965 15486 2991
rect 15653 2965 15683 2991
rect 15752 2965 15782 2991
rect 15838 2965 15868 2991
rect 15922 2965 15952 2991
rect 16030 2965 16060 2991
rect 16114 2965 16144 2991
rect 16278 2965 16308 2991
rect 16497 2965 16527 2991
rect 16594 2965 16624 2991
rect 14677 2816 14707 2831
rect 14644 2786 14707 2816
rect 14644 2733 14674 2786
rect 14761 2742 14791 2831
rect 15028 2794 15058 2881
rect 15120 2843 15150 2881
rect 14620 2717 14674 2733
rect 14620 2683 14630 2717
rect 14664 2683 14674 2717
rect 14716 2732 14791 2742
rect 14716 2698 14732 2732
rect 14766 2698 14791 2732
rect 14929 2778 15058 2794
rect 15104 2833 15170 2843
rect 15104 2799 15120 2833
rect 15154 2799 15170 2833
rect 15104 2789 15170 2799
rect 14929 2744 14939 2778
rect 14973 2764 15058 2778
rect 14973 2744 15046 2764
rect 15219 2747 15249 2881
rect 15359 2823 15389 2881
rect 15359 2807 15414 2823
rect 15359 2773 15369 2807
rect 15403 2773 15414 2807
rect 15359 2757 15414 2773
rect 14929 2728 15046 2744
rect 14716 2688 14791 2698
rect 14620 2667 14674 2683
rect 14644 2644 14674 2667
rect 14644 2614 14707 2644
rect 14677 2599 14707 2614
rect 14761 2599 14791 2688
rect 15016 2599 15046 2728
rect 15111 2717 15249 2747
rect 15111 2687 15142 2717
rect 15088 2671 15142 2687
rect 15088 2637 15098 2671
rect 15132 2637 15142 2671
rect 15088 2621 15142 2637
rect 15184 2665 15250 2675
rect 15184 2631 15200 2665
rect 15234 2631 15250 2665
rect 15184 2621 15250 2631
rect 15111 2587 15141 2621
rect 15207 2587 15237 2621
rect 15373 2599 15403 2757
rect 15456 2687 15486 2881
rect 15653 2782 15683 2797
rect 15577 2752 15683 2782
rect 15577 2735 15607 2752
rect 15541 2719 15607 2735
rect 15445 2671 15499 2687
rect 15445 2637 15455 2671
rect 15489 2637 15499 2671
rect 15541 2685 15551 2719
rect 15585 2685 15607 2719
rect 15752 2747 15782 2881
rect 15838 2849 15868 2881
rect 15824 2833 15878 2849
rect 15824 2799 15834 2833
rect 15868 2799 15878 2833
rect 15824 2783 15878 2799
rect 15752 2735 15802 2747
rect 15752 2723 15815 2735
rect 15752 2717 15839 2723
rect 15773 2707 15839 2717
rect 15773 2705 15795 2707
rect 15541 2669 15607 2685
rect 15577 2643 15607 2669
rect 15676 2659 15743 2675
rect 15445 2621 15499 2637
rect 15445 2599 15475 2621
rect 15676 2625 15699 2659
rect 15733 2625 15743 2659
rect 15676 2609 15743 2625
rect 15785 2673 15795 2705
rect 15829 2673 15839 2707
rect 15785 2657 15839 2673
rect 15922 2697 15952 2881
rect 16030 2725 16060 2881
rect 16114 2833 16144 2881
rect 16102 2817 16156 2833
rect 16102 2783 16112 2817
rect 16146 2783 16156 2817
rect 16102 2767 16156 2783
rect 16025 2709 16079 2725
rect 15922 2681 15983 2697
rect 15922 2661 15939 2681
rect 15676 2587 15706 2609
rect 15785 2587 15815 2657
rect 15881 2647 15939 2661
rect 15973 2647 15983 2681
rect 16025 2675 16035 2709
rect 16069 2675 16079 2709
rect 16025 2659 16079 2675
rect 15881 2631 15983 2647
rect 15881 2599 15911 2631
rect 16030 2599 16060 2659
rect 16121 2599 16151 2767
rect 16497 2801 16527 2837
rect 16486 2771 16527 2801
rect 16278 2733 16308 2765
rect 16486 2733 16516 2771
rect 16594 2733 16624 2765
rect 16207 2717 16516 2733
rect 16207 2683 16235 2717
rect 16269 2683 16516 2717
rect 16207 2667 16516 2683
rect 16565 2717 16624 2733
rect 16565 2683 16575 2717
rect 16609 2683 16624 2717
rect 16565 2667 16624 2683
rect 16309 2645 16339 2667
rect 16486 2644 16516 2667
rect 16594 2645 16624 2667
rect 17192 3494 17258 3510
rect 17192 3460 17208 3494
rect 17242 3460 17258 3494
rect 17192 3444 17258 3460
rect 17210 3413 17240 3444
rect 17210 2782 17240 2813
rect 17192 2766 17258 2782
rect 17192 2732 17208 2766
rect 17242 2732 17258 2766
rect 17192 2716 17258 2732
rect 16486 2614 16527 2644
rect 16497 2599 16527 2614
rect 14677 2489 14707 2515
rect 14761 2489 14791 2515
rect 15016 2489 15046 2515
rect 15111 2489 15141 2515
rect 15207 2489 15237 2515
rect 15373 2489 15403 2515
rect 15445 2489 15475 2515
rect 15577 2489 15607 2515
rect 15676 2489 15706 2515
rect 15785 2489 15815 2515
rect 15881 2489 15911 2515
rect 16030 2489 16060 2515
rect 16121 2489 16151 2515
rect 16309 2489 16339 2515
rect 16497 2489 16527 2515
rect 16594 2489 16624 2515
rect 17192 2406 17258 2422
rect 17192 2372 17208 2406
rect 17242 2372 17258 2406
rect 17192 2356 17258 2372
rect 17210 2334 17240 2356
rect 17210 2112 17240 2134
rect 218 1944 418 1960
rect 218 1910 234 1944
rect 402 1910 418 1944
rect 218 1872 418 1910
rect 598 1944 798 1960
rect 598 1910 614 1944
rect 782 1910 798 1944
rect 598 1872 798 1910
rect 978 1944 1178 1960
rect 978 1910 994 1944
rect 1162 1910 1178 1944
rect 978 1872 1178 1910
rect 1358 1944 1558 1960
rect 1358 1910 1374 1944
rect 1542 1910 1558 1944
rect 1358 1872 1558 1910
rect 1738 1944 1938 1960
rect 1738 1910 1754 1944
rect 1922 1910 1938 1944
rect 1738 1872 1938 1910
rect 2118 1944 2318 1960
rect 2118 1910 2134 1944
rect 2302 1910 2318 1944
rect 2118 1872 2318 1910
rect 2498 1944 2698 1960
rect 2498 1910 2514 1944
rect 2682 1910 2698 1944
rect 2498 1872 2698 1910
rect 2878 1944 3078 1960
rect 2878 1910 2894 1944
rect 3062 1910 3078 1944
rect 2878 1872 3078 1910
rect 17192 2096 17258 2112
rect 17192 2062 17208 2096
rect 17242 2062 17258 2096
rect 17192 2046 17258 2062
rect 218 1634 418 1672
rect 218 1600 234 1634
rect 402 1600 418 1634
rect 218 1584 418 1600
rect 598 1634 798 1672
rect 598 1600 614 1634
rect 782 1600 798 1634
rect 598 1584 798 1600
rect 978 1634 1178 1672
rect 978 1600 994 1634
rect 1162 1600 1178 1634
rect 978 1584 1178 1600
rect 1358 1634 1558 1672
rect 1358 1600 1374 1634
rect 1542 1600 1558 1634
rect 1358 1584 1558 1600
rect 1738 1634 1938 1672
rect 1738 1600 1754 1634
rect 1922 1600 1938 1634
rect 1738 1584 1938 1600
rect 2118 1634 2318 1672
rect 2118 1600 2134 1634
rect 2302 1600 2318 1634
rect 2118 1584 2318 1600
rect 2498 1634 2698 1672
rect 2498 1600 2514 1634
rect 2682 1600 2698 1634
rect 2498 1584 2698 1600
rect 2878 1634 3078 1672
rect 2878 1600 2894 1634
rect 3062 1600 3078 1634
rect 2878 1584 3078 1600
rect 218 1526 418 1542
rect 218 1492 234 1526
rect 402 1492 418 1526
rect 218 1454 418 1492
rect 598 1526 798 1542
rect 598 1492 614 1526
rect 782 1492 798 1526
rect 598 1454 798 1492
rect 978 1526 1178 1542
rect 978 1492 994 1526
rect 1162 1492 1178 1526
rect 978 1454 1178 1492
rect 1358 1526 1558 1542
rect 1358 1492 1374 1526
rect 1542 1492 1558 1526
rect 1358 1454 1558 1492
rect 1738 1526 1938 1542
rect 1738 1492 1754 1526
rect 1922 1492 1938 1526
rect 1738 1454 1938 1492
rect 2118 1526 2318 1542
rect 2118 1492 2134 1526
rect 2302 1492 2318 1526
rect 2118 1454 2318 1492
rect 2498 1526 2698 1542
rect 2498 1492 2514 1526
rect 2682 1492 2698 1526
rect 2498 1454 2698 1492
rect 2878 1526 3078 1542
rect 2878 1492 2894 1526
rect 3062 1492 3078 1526
rect 2878 1454 3078 1492
rect 218 1216 418 1254
rect 218 1182 234 1216
rect 402 1182 418 1216
rect 218 1166 418 1182
rect 598 1216 798 1254
rect 598 1182 614 1216
rect 782 1182 798 1216
rect 598 1166 798 1182
rect 978 1216 1178 1254
rect 978 1182 994 1216
rect 1162 1182 1178 1216
rect 978 1166 1178 1182
rect 1358 1216 1558 1254
rect 1358 1182 1374 1216
rect 1542 1182 1558 1216
rect 1358 1166 1558 1182
rect 1738 1216 1938 1254
rect 1738 1182 1754 1216
rect 1922 1182 1938 1216
rect 1738 1166 1938 1182
rect 2118 1216 2318 1254
rect 2118 1182 2134 1216
rect 2302 1182 2318 1216
rect 2118 1166 2318 1182
rect 2498 1216 2698 1254
rect 2498 1182 2514 1216
rect 2682 1182 2698 1216
rect 2498 1166 2698 1182
rect 2878 1216 3078 1254
rect 2878 1182 2894 1216
rect 3062 1182 3078 1216
rect 2878 1166 3078 1182
rect 218 1108 418 1124
rect 218 1074 234 1108
rect 402 1074 418 1108
rect 218 1036 418 1074
rect 598 1108 798 1124
rect 598 1074 614 1108
rect 782 1074 798 1108
rect 598 1036 798 1074
rect 978 1108 1178 1124
rect 978 1074 994 1108
rect 1162 1074 1178 1108
rect 978 1036 1178 1074
rect 1358 1108 1558 1124
rect 1358 1074 1374 1108
rect 1542 1074 1558 1108
rect 1358 1036 1558 1074
rect 1738 1108 1938 1124
rect 1738 1074 1754 1108
rect 1922 1074 1938 1108
rect 1738 1036 1938 1074
rect 2118 1108 2318 1124
rect 2118 1074 2134 1108
rect 2302 1074 2318 1108
rect 2118 1036 2318 1074
rect 2498 1108 2698 1124
rect 2498 1074 2514 1108
rect 2682 1074 2698 1108
rect 2498 1036 2698 1074
rect 2878 1108 3078 1124
rect 2878 1074 2894 1108
rect 3062 1074 3078 1108
rect 2878 1036 3078 1074
rect 218 798 418 836
rect 218 764 234 798
rect 402 764 418 798
rect 218 748 418 764
rect 598 798 798 836
rect 598 764 614 798
rect 782 764 798 798
rect 598 748 798 764
rect 978 798 1178 836
rect 978 764 994 798
rect 1162 764 1178 798
rect 978 748 1178 764
rect 1358 798 1558 836
rect 1358 764 1374 798
rect 1542 764 1558 798
rect 1358 748 1558 764
rect 1738 798 1938 836
rect 1738 764 1754 798
rect 1922 764 1938 798
rect 1738 748 1938 764
rect 2118 798 2318 836
rect 2118 764 2134 798
rect 2302 764 2318 798
rect 2118 748 2318 764
rect 2498 798 2698 836
rect 2498 764 2514 798
rect 2682 764 2698 798
rect 2498 748 2698 764
rect 2878 798 3078 836
rect 2878 764 2894 798
rect 3062 764 3078 798
rect 2878 748 3078 764
rect 218 690 418 706
rect 218 656 234 690
rect 402 656 418 690
rect 218 618 418 656
rect 598 690 798 706
rect 598 656 614 690
rect 782 656 798 690
rect 598 618 798 656
rect 978 690 1178 706
rect 978 656 994 690
rect 1162 656 1178 690
rect 978 618 1178 656
rect 1358 690 1558 706
rect 1358 656 1374 690
rect 1542 656 1558 690
rect 1358 618 1558 656
rect 1738 690 1938 706
rect 1738 656 1754 690
rect 1922 656 1938 690
rect 1738 618 1938 656
rect 2118 690 2318 706
rect 2118 656 2134 690
rect 2302 656 2318 690
rect 2118 618 2318 656
rect 2498 690 2698 706
rect 2498 656 2514 690
rect 2682 656 2698 690
rect 2498 618 2698 656
rect 2878 690 3078 706
rect 2878 656 2894 690
rect 3062 656 3078 690
rect 2878 618 3078 656
rect 218 380 418 418
rect 218 346 234 380
rect 402 346 418 380
rect 218 330 418 346
rect 598 380 798 418
rect 598 346 614 380
rect 782 346 798 380
rect 598 330 798 346
rect 978 380 1178 418
rect 978 346 994 380
rect 1162 346 1178 380
rect 978 330 1178 346
rect 1358 380 1558 418
rect 1358 346 1374 380
rect 1542 346 1558 380
rect 1358 330 1558 346
rect 1738 380 1938 418
rect 1738 346 1754 380
rect 1922 346 1938 380
rect 1738 330 1938 346
rect 2118 380 2318 418
rect 2118 346 2134 380
rect 2302 346 2318 380
rect 2118 330 2318 346
rect 2498 380 2698 418
rect 2498 346 2514 380
rect 2682 346 2698 380
rect 2498 330 2698 346
rect 2878 380 3078 418
rect 2878 346 2894 380
rect 3062 346 3078 380
rect 2878 330 3078 346
<< polycont >>
rect 874 10988 908 11022
rect 874 10478 908 10512
rect 5870 6047 6038 6081
rect 6128 6047 6296 6081
rect 6386 6047 6554 6081
rect 6644 6047 6812 6081
rect 6902 6047 7070 6081
rect 7160 6047 7328 6081
rect 7530 6047 7698 6081
rect 7910 6047 8078 6081
rect 8168 6047 8336 6081
rect 8426 6047 8594 6081
rect 8684 6047 8852 6081
rect 8942 6047 9110 6081
rect 9330 6047 9498 6081
rect 9588 6047 9756 6081
rect 9846 6047 10014 6081
rect 10104 6047 10272 6081
rect 10362 6047 10530 6081
rect 10750 6047 10918 6081
rect 11130 6047 11298 6081
rect 11388 6047 11556 6081
rect 11646 6047 11814 6081
rect 11904 6047 12072 6081
rect 12162 6047 12330 6081
rect 12420 6047 12588 6081
rect 5870 5719 6038 5753
rect 6128 5719 6296 5753
rect 6386 5719 6554 5753
rect 6644 5719 6812 5753
rect 6902 5719 7070 5753
rect 7160 5719 7328 5753
rect 7530 5719 7698 5753
rect 7910 5719 8078 5753
rect 8168 5719 8336 5753
rect 8426 5719 8594 5753
rect 8684 5719 8852 5753
rect 8942 5719 9110 5753
rect 9330 5719 9498 5753
rect 9588 5719 9756 5753
rect 9846 5719 10014 5753
rect 10104 5719 10272 5753
rect 10362 5719 10530 5753
rect 10750 5719 10918 5753
rect 11130 5719 11298 5753
rect 11388 5719 11556 5753
rect 11646 5719 11814 5753
rect 11904 5719 12072 5753
rect 12162 5719 12330 5753
rect 12420 5719 12588 5753
rect 1830 5027 1998 5061
rect 2210 5027 2378 5061
rect 2590 5027 3558 5061
rect 3770 5027 3938 5061
rect 1830 4499 1998 4533
rect 2210 4499 2378 4533
rect 2590 4499 3558 4533
rect 3770 4499 3938 4533
rect 450 4347 618 4381
rect 830 4347 998 4381
rect 1088 4347 1256 4381
rect 1470 4347 1638 4381
rect 1728 4347 1896 4381
rect 1986 4347 2154 4381
rect 2244 4347 2412 4381
rect 2630 4347 2798 4381
rect 2888 4347 3056 4381
rect 3146 4347 3314 4381
rect 3404 4347 3572 4381
rect 3790 4347 3958 4381
rect 450 3819 618 3853
rect 830 3819 998 3853
rect 1088 3819 1256 3853
rect 1470 3819 1638 3853
rect 1728 3819 1896 3853
rect 1986 3819 2154 3853
rect 2244 3819 2412 3853
rect 2630 3819 2798 3853
rect 2888 3819 3056 3853
rect 3146 3819 3314 3853
rect 3404 3819 3572 3853
rect 3790 3819 3958 3853
rect 5900 5120 6068 5154
rect 6158 5120 6326 5154
rect 6416 5120 6584 5154
rect 6674 5120 6842 5154
rect 6932 5120 7100 5154
rect 7190 5120 7358 5154
rect 7448 5120 7616 5154
rect 7706 5120 7874 5154
rect 7964 5120 8132 5154
rect 8222 5120 8390 5154
rect 8480 5120 8648 5154
rect 8738 5120 8906 5154
rect 8996 5120 9164 5154
rect 9254 5120 9422 5154
rect 9512 5120 9680 5154
rect 9770 5120 9938 5154
rect 10028 5120 10196 5154
rect 10286 5120 10454 5154
rect 10544 5120 10712 5154
rect 10802 5120 10970 5154
rect 11060 5120 11228 5154
rect 11318 5120 11486 5154
rect 5900 4810 6068 4844
rect 6158 4810 6326 4844
rect 6416 4810 6584 4844
rect 6674 4810 6842 4844
rect 6932 4810 7100 4844
rect 7190 4810 7358 4844
rect 7448 4810 7616 4844
rect 7706 4810 7874 4844
rect 7964 4810 8132 4844
rect 8222 4810 8390 4844
rect 8480 4810 8648 4844
rect 8738 4810 8906 4844
rect 8996 4810 9164 4844
rect 9254 4810 9422 4844
rect 9512 4810 9680 4844
rect 9770 4810 9938 4844
rect 10028 4810 10196 4844
rect 10286 4810 10454 4844
rect 10544 4810 10712 4844
rect 10802 4810 10970 4844
rect 11060 4810 11228 4844
rect 11318 4810 11486 4844
rect 5994 4286 6162 4320
rect 6252 4286 6420 4320
rect 6510 4286 6678 4320
rect 6914 4286 7082 4320
rect 7172 4286 7340 4320
rect 7430 4286 7598 4320
rect 7688 4286 7856 4320
rect 7946 4286 8114 4320
rect 8204 4286 8372 4320
rect 8462 4286 8630 4320
rect 8720 4286 8888 4320
rect 8978 4286 9146 4320
rect 9236 4286 9404 4320
rect 9494 4286 9662 4320
rect 9752 4286 9920 4320
rect 10010 4286 10178 4320
rect 10268 4286 10436 4320
rect 10526 4286 10694 4320
rect 10784 4286 10952 4320
rect 11042 4286 11210 4320
rect 11300 4286 11468 4320
rect 11558 4286 11726 4320
rect 11816 4286 11984 4320
rect 12074 4286 12242 4320
rect 5994 3976 6162 4010
rect 6252 3976 6420 4010
rect 6510 3976 6678 4010
rect 6914 3976 7082 4010
rect 7172 3976 7340 4010
rect 7430 3976 7598 4010
rect 7688 3976 7856 4010
rect 7946 3976 8114 4010
rect 8204 3976 8372 4010
rect 8462 3976 8630 4010
rect 8720 3976 8888 4010
rect 8978 3976 9146 4010
rect 9236 3976 9404 4010
rect 9494 3976 9662 4010
rect 9752 3976 9920 4010
rect 10010 3976 10178 4010
rect 10268 3976 10436 4010
rect 10526 3976 10694 4010
rect 10784 3976 10952 4010
rect 11042 3976 11210 4010
rect 11300 3976 11468 4010
rect 11558 3976 11726 4010
rect 11816 3976 11984 4010
rect 12074 3976 12242 4010
rect 430 3107 598 3141
rect 810 3107 978 3141
rect 1068 3107 1236 3141
rect 1326 3107 1494 3141
rect 1584 3107 1752 3141
rect 1842 3107 2010 3141
rect 2100 3107 2268 3141
rect 2358 3107 2526 3141
rect 2616 3107 2784 3141
rect 2990 3107 3158 3141
rect 430 2579 598 2613
rect 810 2579 978 2613
rect 1068 2579 1236 2613
rect 1326 2579 1494 2613
rect 1584 2579 1752 2613
rect 1842 2579 2010 2613
rect 2100 2579 2268 2613
rect 2358 2579 2526 2613
rect 2616 2579 2784 2613
rect 2990 2579 3158 2613
rect 14630 2683 14664 2717
rect 14732 2698 14766 2732
rect 15120 2799 15154 2833
rect 14939 2744 14973 2778
rect 15369 2773 15403 2807
rect 15098 2637 15132 2671
rect 15200 2631 15234 2665
rect 15455 2637 15489 2671
rect 15551 2685 15585 2719
rect 15834 2799 15868 2833
rect 15699 2625 15733 2659
rect 15795 2673 15829 2707
rect 16112 2783 16146 2817
rect 15939 2647 15973 2681
rect 16035 2675 16069 2709
rect 16235 2683 16269 2717
rect 16575 2683 16609 2717
rect 17208 3460 17242 3494
rect 17208 2732 17242 2766
rect 17208 2372 17242 2406
rect 234 1910 402 1944
rect 614 1910 782 1944
rect 994 1910 1162 1944
rect 1374 1910 1542 1944
rect 1754 1910 1922 1944
rect 2134 1910 2302 1944
rect 2514 1910 2682 1944
rect 2894 1910 3062 1944
rect 17208 2062 17242 2096
rect 234 1600 402 1634
rect 614 1600 782 1634
rect 994 1600 1162 1634
rect 1374 1600 1542 1634
rect 1754 1600 1922 1634
rect 2134 1600 2302 1634
rect 2514 1600 2682 1634
rect 2894 1600 3062 1634
rect 234 1492 402 1526
rect 614 1492 782 1526
rect 994 1492 1162 1526
rect 1374 1492 1542 1526
rect 1754 1492 1922 1526
rect 2134 1492 2302 1526
rect 2514 1492 2682 1526
rect 2894 1492 3062 1526
rect 234 1182 402 1216
rect 614 1182 782 1216
rect 994 1182 1162 1216
rect 1374 1182 1542 1216
rect 1754 1182 1922 1216
rect 2134 1182 2302 1216
rect 2514 1182 2682 1216
rect 2894 1182 3062 1216
rect 234 1074 402 1108
rect 614 1074 782 1108
rect 994 1074 1162 1108
rect 1374 1074 1542 1108
rect 1754 1074 1922 1108
rect 2134 1074 2302 1108
rect 2514 1074 2682 1108
rect 2894 1074 3062 1108
rect 234 764 402 798
rect 614 764 782 798
rect 994 764 1162 798
rect 1374 764 1542 798
rect 1754 764 1922 798
rect 2134 764 2302 798
rect 2514 764 2682 798
rect 2894 764 3062 798
rect 234 656 402 690
rect 614 656 782 690
rect 994 656 1162 690
rect 1374 656 1542 690
rect 1754 656 1922 690
rect 2134 656 2302 690
rect 2514 656 2682 690
rect 2894 656 3062 690
rect 234 346 402 380
rect 614 346 782 380
rect 994 346 1162 380
rect 1374 346 1542 380
rect 1754 346 1922 380
rect 2134 346 2302 380
rect 2514 346 2682 380
rect 2894 346 3062 380
<< xpolycontact >>
rect 6126 30818 6196 31250
rect 6126 29386 6196 29818
rect 14550 5320 14620 5752
rect 14550 3988 14620 4420
rect 14716 5320 14786 5752
rect 14716 3988 14786 4420
rect 14882 5320 14952 5752
rect 14882 3988 14952 4420
rect 15048 5320 15118 5752
rect 15048 3988 15118 4420
rect 15214 5320 15284 5752
rect 15214 3988 15284 4420
rect 15380 5320 15450 5752
rect 15380 3988 15450 4420
rect 15546 5320 15616 5752
rect 15546 3988 15616 4420
rect 15712 5320 15782 5752
rect 15712 3988 15782 4420
rect 16024 5320 16094 5752
rect 16024 3988 16094 4420
rect 16190 5320 16260 5752
rect 16190 3988 16260 4420
rect 16356 5320 16426 5752
rect 16356 3988 16426 4420
rect 16522 5320 16592 5752
rect 16522 3988 16592 4420
rect 16688 5320 16758 5752
rect 16688 3988 16758 4420
rect 16854 5320 16924 5752
rect 16854 3988 16924 4420
rect 17020 5320 17090 5752
rect 17020 3988 17090 4420
rect 17186 5320 17256 5752
rect 17186 3988 17256 4420
<< xpolyres >>
rect 6126 29818 6196 30818
rect 14550 4420 14620 5320
rect 14716 4420 14786 5320
rect 14882 4420 14952 5320
rect 15048 4420 15118 5320
rect 15214 4420 15284 5320
rect 15380 4420 15450 5320
rect 15546 4420 15616 5320
rect 15712 4420 15782 5320
rect 16024 4420 16094 5320
rect 16190 4420 16260 5320
rect 16356 4420 16426 5320
rect 16522 4420 16592 5320
rect 16688 4420 16758 5320
rect 16854 4420 16924 5320
rect 17020 4420 17090 5320
rect 17186 4420 17256 5320
<< locali >>
rect 5996 31346 6092 31380
rect 6230 31346 6326 31380
rect 5996 31284 6030 31346
rect 6292 31284 6326 31346
rect 5996 29290 6030 29352
rect 6292 29290 6326 29352
rect 5996 29256 6092 29290
rect 6230 29256 6326 29290
rect 716 11090 812 11124
rect 970 11090 1066 11124
rect 716 11028 750 11090
rect 1032 11028 1066 11090
rect 858 10988 874 11022
rect 908 10988 924 11022
rect 830 10938 864 10954
rect 830 10546 864 10562
rect 918 10938 952 10954
rect 918 10546 952 10562
rect 858 10478 874 10512
rect 908 10478 924 10512
rect 716 10410 750 10472
rect 1032 10410 1066 10472
rect 716 10376 812 10410
rect 970 10376 1066 10410
rect 5683 6183 5743 6217
rect 12717 6183 12777 6217
rect 5683 6157 5717 6183
rect 12743 6157 12777 6183
rect 5854 6047 5870 6081
rect 6038 6047 6054 6081
rect 6112 6047 6128 6081
rect 6296 6047 6312 6081
rect 6370 6047 6386 6081
rect 6554 6047 6570 6081
rect 6628 6047 6644 6081
rect 6812 6047 6828 6081
rect 6886 6047 6902 6081
rect 7070 6047 7086 6081
rect 7144 6047 7160 6081
rect 7328 6047 7344 6081
rect 7514 6047 7530 6081
rect 7698 6047 7714 6081
rect 7894 6047 7910 6081
rect 8078 6047 8094 6081
rect 8152 6047 8168 6081
rect 8336 6047 8352 6081
rect 8410 6047 8426 6081
rect 8594 6047 8610 6081
rect 8668 6047 8684 6081
rect 8852 6047 8868 6081
rect 8926 6047 8942 6081
rect 9110 6047 9126 6081
rect 9314 6047 9330 6081
rect 9498 6047 9514 6081
rect 9572 6047 9588 6081
rect 9756 6047 9772 6081
rect 9830 6047 9846 6081
rect 10014 6047 10030 6081
rect 10088 6047 10104 6081
rect 10272 6047 10288 6081
rect 10346 6047 10362 6081
rect 10530 6047 10546 6081
rect 10734 6047 10750 6081
rect 10918 6047 10934 6081
rect 11114 6047 11130 6081
rect 11298 6047 11314 6081
rect 11372 6047 11388 6081
rect 11556 6047 11572 6081
rect 11630 6047 11646 6081
rect 11814 6047 11830 6081
rect 11888 6047 11904 6081
rect 12072 6047 12088 6081
rect 12146 6047 12162 6081
rect 12330 6047 12346 6081
rect 12404 6047 12420 6081
rect 12588 6047 12604 6081
rect 5808 5988 5842 6004
rect 5808 5796 5842 5812
rect 6066 5988 6100 6004
rect 6066 5796 6100 5812
rect 6324 5988 6358 6004
rect 6324 5796 6358 5812
rect 6582 5988 6616 6004
rect 6582 5796 6616 5812
rect 6840 5988 6874 6004
rect 6840 5796 6874 5812
rect 7098 5988 7132 6004
rect 7098 5796 7132 5812
rect 7356 5988 7390 6004
rect 7356 5796 7390 5812
rect 7468 5988 7502 6004
rect 7468 5796 7502 5812
rect 7726 5988 7760 6004
rect 7726 5796 7760 5812
rect 7848 5988 7882 6004
rect 7848 5796 7882 5812
rect 8106 5988 8140 6004
rect 8106 5796 8140 5812
rect 8364 5988 8398 6004
rect 8364 5796 8398 5812
rect 8622 5988 8656 6004
rect 8622 5796 8656 5812
rect 8880 5988 8914 6004
rect 8880 5796 8914 5812
rect 9138 5988 9172 6004
rect 9138 5796 9172 5812
rect 9268 5988 9302 6004
rect 9268 5796 9302 5812
rect 9526 5988 9560 6004
rect 9526 5796 9560 5812
rect 9784 5988 9818 6004
rect 9784 5796 9818 5812
rect 10042 5988 10076 6004
rect 10042 5796 10076 5812
rect 10300 5988 10334 6004
rect 10300 5796 10334 5812
rect 10558 5988 10592 6004
rect 10558 5796 10592 5812
rect 10688 5988 10722 6004
rect 10688 5796 10722 5812
rect 10946 5988 10980 6004
rect 10946 5796 10980 5812
rect 11068 5988 11102 6004
rect 11068 5796 11102 5812
rect 11326 5988 11360 6004
rect 11326 5796 11360 5812
rect 11584 5988 11618 6004
rect 11584 5796 11618 5812
rect 11842 5988 11876 6004
rect 11842 5796 11876 5812
rect 12100 5988 12134 6004
rect 12100 5796 12134 5812
rect 12358 5988 12392 6004
rect 12358 5796 12392 5812
rect 12616 5988 12650 6004
rect 12616 5796 12650 5812
rect 5854 5719 5870 5753
rect 6038 5719 6054 5753
rect 6112 5719 6128 5753
rect 6296 5719 6312 5753
rect 6370 5719 6386 5753
rect 6554 5719 6570 5753
rect 6628 5719 6644 5753
rect 6812 5719 6828 5753
rect 6886 5719 6902 5753
rect 7070 5719 7086 5753
rect 7144 5719 7160 5753
rect 7328 5719 7344 5753
rect 7514 5719 7530 5753
rect 7698 5719 7714 5753
rect 7894 5719 7910 5753
rect 8078 5719 8094 5753
rect 8152 5719 8168 5753
rect 8336 5719 8352 5753
rect 8410 5719 8426 5753
rect 8594 5719 8610 5753
rect 8668 5719 8684 5753
rect 8852 5719 8868 5753
rect 8926 5719 8942 5753
rect 9110 5719 9126 5753
rect 9314 5719 9330 5753
rect 9498 5719 9514 5753
rect 9572 5719 9588 5753
rect 9756 5719 9772 5753
rect 9830 5719 9846 5753
rect 10014 5719 10030 5753
rect 10088 5719 10104 5753
rect 10272 5719 10288 5753
rect 10346 5719 10362 5753
rect 10530 5719 10546 5753
rect 10734 5719 10750 5753
rect 10918 5719 10934 5753
rect 11114 5719 11130 5753
rect 11298 5719 11314 5753
rect 11372 5719 11388 5753
rect 11556 5719 11572 5753
rect 11630 5719 11646 5753
rect 11814 5719 11830 5753
rect 11888 5719 11904 5753
rect 12072 5719 12088 5753
rect 12146 5719 12162 5753
rect 12330 5719 12346 5753
rect 12404 5719 12420 5753
rect 12588 5719 12604 5753
rect 5683 5637 5717 5663
rect 12743 5637 12777 5663
rect 5683 5603 5743 5637
rect 12717 5603 12777 5637
rect 243 5223 303 5257
rect 4137 5223 4197 5257
rect 243 5197 277 5223
rect 4163 5197 4197 5223
rect 1814 5027 1830 5061
rect 1998 5027 2014 5061
rect 2194 5027 2210 5061
rect 2378 5027 2394 5061
rect 2574 5027 2590 5061
rect 3558 5027 3574 5061
rect 3754 5027 3770 5061
rect 3938 5027 3954 5061
rect 1768 4968 1802 4984
rect 1768 4576 1802 4592
rect 2026 4968 2060 4984
rect 2026 4576 2060 4592
rect 2148 4968 2182 4984
rect 2148 4576 2182 4592
rect 2406 4968 2440 4984
rect 2406 4576 2440 4592
rect 2528 4968 2562 4984
rect 2528 4576 2562 4592
rect 3586 4968 3620 4984
rect 3586 4576 3620 4592
rect 3708 4968 3742 4984
rect 3708 4576 3742 4592
rect 3966 4968 4000 4984
rect 3966 4576 4000 4592
rect 1814 4499 1830 4533
rect 1998 4499 2014 4533
rect 2194 4499 2210 4533
rect 2378 4499 2394 4533
rect 2574 4499 2590 4533
rect 3558 4499 3574 4533
rect 3754 4499 3770 4533
rect 3938 4499 3954 4533
rect 434 4347 450 4381
rect 618 4347 634 4381
rect 814 4347 830 4381
rect 998 4347 1014 4381
rect 1072 4347 1088 4381
rect 1256 4347 1272 4381
rect 1454 4347 1470 4381
rect 1638 4347 1654 4381
rect 1712 4347 1728 4381
rect 1896 4347 1912 4381
rect 1970 4347 1986 4381
rect 2154 4347 2170 4381
rect 2228 4347 2244 4381
rect 2412 4347 2428 4381
rect 2614 4347 2630 4381
rect 2798 4347 2814 4381
rect 2872 4347 2888 4381
rect 3056 4347 3072 4381
rect 3130 4347 3146 4381
rect 3314 4347 3330 4381
rect 3388 4347 3404 4381
rect 3572 4347 3588 4381
rect 3774 4347 3790 4381
rect 3958 4347 3974 4381
rect 388 4288 422 4304
rect 388 3896 422 3912
rect 646 4288 680 4304
rect 646 3896 680 3912
rect 768 4288 802 4304
rect 768 3896 802 3912
rect 1026 4288 1060 4304
rect 1026 3896 1060 3912
rect 1284 4288 1318 4304
rect 1284 3896 1318 3912
rect 1408 4288 1442 4304
rect 1408 3896 1442 3912
rect 1666 4288 1700 4304
rect 1666 3896 1700 3912
rect 1924 4288 1958 4304
rect 1924 3896 1958 3912
rect 2182 4288 2216 4304
rect 2182 3896 2216 3912
rect 2440 4288 2474 4304
rect 2440 3896 2474 3912
rect 2568 4288 2602 4304
rect 2568 3896 2602 3912
rect 2826 4288 2860 4304
rect 2826 3896 2860 3912
rect 3084 4288 3118 4304
rect 3084 3896 3118 3912
rect 3342 4288 3376 4304
rect 3342 3896 3376 3912
rect 3600 4288 3634 4304
rect 3600 3896 3634 3912
rect 3728 4288 3762 4304
rect 3728 3896 3762 3912
rect 3986 4288 4020 4304
rect 3986 3896 4020 3912
rect 434 3819 450 3853
rect 618 3819 634 3853
rect 814 3819 830 3853
rect 998 3819 1014 3853
rect 1072 3819 1088 3853
rect 1256 3819 1272 3853
rect 1454 3819 1470 3853
rect 1638 3819 1654 3853
rect 1712 3819 1728 3853
rect 1896 3819 1912 3853
rect 1970 3819 1986 3853
rect 2154 3819 2170 3853
rect 2228 3819 2244 3853
rect 2412 3819 2428 3853
rect 2614 3819 2630 3853
rect 2798 3819 2814 3853
rect 2872 3819 2888 3853
rect 3056 3819 3072 3853
rect 3130 3819 3146 3853
rect 3314 3819 3330 3853
rect 3388 3819 3404 3853
rect 3572 3819 3588 3853
rect 3774 3819 3790 3853
rect 3958 3819 3974 3853
rect 243 3697 277 3723
rect 5736 5230 5832 5264
rect 11960 5230 12056 5264
rect 5736 5168 5770 5230
rect 12022 5168 12056 5230
rect 5884 5120 5900 5154
rect 6068 5120 6084 5154
rect 6142 5120 6158 5154
rect 6326 5120 6342 5154
rect 6400 5120 6416 5154
rect 6584 5120 6600 5154
rect 6658 5120 6674 5154
rect 6842 5120 6858 5154
rect 6916 5120 6932 5154
rect 7100 5120 7116 5154
rect 7174 5120 7180 5154
rect 7358 5120 7374 5154
rect 7432 5120 7448 5154
rect 7616 5120 7632 5154
rect 7690 5120 7706 5154
rect 7874 5120 7890 5154
rect 7948 5120 7960 5154
rect 8132 5120 8148 5154
rect 8206 5120 8220 5154
rect 8390 5120 8406 5154
rect 8464 5120 8480 5154
rect 8648 5120 8664 5154
rect 8722 5120 8738 5154
rect 8906 5120 8922 5154
rect 8980 5120 8996 5154
rect 9164 5120 9180 5154
rect 9238 5120 9254 5154
rect 9422 5120 9438 5154
rect 9496 5120 9512 5154
rect 9680 5120 9696 5154
rect 9754 5120 9770 5154
rect 9938 5120 9954 5154
rect 10012 5120 10020 5154
rect 10196 5120 10212 5154
rect 10270 5120 10280 5154
rect 10454 5120 10470 5154
rect 10528 5120 10544 5154
rect 10712 5120 10728 5154
rect 10786 5120 10802 5154
rect 10970 5120 10986 5154
rect 11044 5120 11060 5154
rect 11228 5120 11244 5154
rect 11302 5120 11318 5154
rect 11486 5120 11502 5154
rect 5838 5070 5872 5086
rect 5838 4878 5872 4894
rect 6096 5070 6130 5086
rect 6096 4878 6130 4894
rect 6354 5070 6388 5086
rect 6354 4878 6388 4894
rect 6612 5070 6646 5086
rect 6612 4878 6646 4894
rect 6870 5070 6904 5086
rect 6870 4878 6904 4894
rect 7128 5070 7162 5086
rect 7128 4878 7162 4894
rect 7386 5070 7420 5086
rect 7386 4878 7420 4894
rect 7644 5070 7678 5086
rect 7644 4878 7678 4894
rect 7902 5070 7936 5086
rect 7902 4878 7936 4894
rect 8160 5070 8194 5086
rect 8160 4878 8194 4894
rect 8418 5070 8452 5086
rect 8418 4878 8452 4894
rect 8676 5070 8710 5086
rect 8676 4878 8710 4894
rect 8934 5070 8968 5086
rect 8934 4878 8968 4894
rect 9192 5070 9226 5086
rect 9192 4878 9226 4894
rect 9450 5070 9484 5086
rect 9450 4878 9484 4894
rect 9708 5070 9742 5086
rect 9708 4878 9742 4894
rect 9966 5070 10000 5086
rect 9966 4878 10000 4894
rect 10224 5070 10258 5086
rect 10224 4878 10258 4894
rect 10482 5070 10516 5086
rect 10482 4878 10516 4894
rect 10740 5070 10774 5086
rect 10740 4878 10774 4894
rect 10998 5070 11032 5086
rect 10998 4878 11032 4894
rect 11256 5070 11290 5086
rect 11256 4878 11290 4894
rect 11514 5070 11548 5086
rect 11514 4878 11548 4894
rect 5736 4750 5770 4812
rect 5884 4810 5900 4844
rect 6068 4810 6084 4844
rect 6142 4810 6158 4844
rect 6326 4810 6342 4844
rect 6400 4810 6416 4844
rect 6584 4810 6600 4844
rect 6658 4810 6674 4844
rect 6842 4810 6858 4844
rect 6916 4810 6932 4844
rect 7100 4810 7116 4844
rect 7174 4810 7190 4844
rect 7358 4810 7374 4844
rect 7432 4840 7448 4844
rect 7432 4810 7440 4840
rect 7616 4810 7632 4844
rect 7690 4840 7706 4844
rect 7690 4810 7700 4840
rect 7874 4810 7890 4844
rect 7948 4810 7964 4844
rect 8132 4810 8148 4844
rect 8206 4810 8222 4844
rect 8390 4810 8406 4844
rect 8464 4810 8480 4844
rect 8648 4810 8664 4844
rect 8722 4810 8738 4844
rect 8906 4810 8922 4844
rect 8980 4810 8996 4844
rect 9164 4810 9180 4844
rect 9238 4810 9254 4844
rect 9422 4810 9438 4844
rect 9496 4810 9512 4844
rect 9680 4810 9696 4844
rect 9754 4840 9770 4844
rect 9754 4810 9760 4840
rect 9938 4810 9954 4844
rect 10012 4810 10028 4844
rect 10196 4810 10212 4844
rect 10270 4810 10286 4844
rect 10454 4810 10470 4844
rect 10528 4840 10544 4844
rect 10528 4810 10540 4840
rect 10712 4810 10728 4844
rect 10786 4840 10802 4844
rect 10786 4810 10800 4840
rect 10970 4810 10986 4844
rect 11044 4810 11060 4844
rect 11228 4810 11244 4844
rect 11302 4810 11318 4844
rect 11486 4810 11502 4844
rect 12022 4750 12056 4812
rect 5736 4716 5832 4750
rect 11960 4716 12056 4750
rect 5816 4390 5912 4424
rect 12440 4390 12536 4424
rect 5816 4328 5850 4390
rect 12502 4328 12536 4390
rect 5978 4286 5994 4320
rect 6162 4286 6178 4320
rect 6236 4286 6252 4320
rect 6420 4286 6436 4320
rect 6494 4286 6510 4320
rect 6678 4286 6694 4320
rect 6898 4286 6914 4320
rect 7082 4286 7098 4320
rect 7156 4286 7172 4320
rect 7340 4286 7356 4320
rect 7414 4286 7430 4320
rect 7598 4286 7614 4320
rect 7672 4286 7688 4320
rect 7856 4286 7872 4320
rect 7930 4286 7946 4320
rect 8114 4286 8130 4320
rect 8188 4286 8204 4320
rect 8372 4286 8388 4320
rect 8446 4286 8462 4320
rect 8630 4286 8646 4320
rect 8704 4286 8720 4320
rect 8888 4286 8904 4320
rect 8962 4286 8978 4320
rect 9146 4286 9162 4320
rect 9220 4286 9236 4320
rect 9404 4286 9420 4320
rect 9478 4286 9494 4320
rect 9662 4286 9678 4320
rect 9736 4286 9752 4320
rect 9920 4286 9936 4320
rect 9994 4286 10010 4320
rect 10178 4286 10194 4320
rect 10252 4286 10268 4320
rect 10436 4286 10452 4320
rect 10510 4286 10526 4320
rect 10694 4286 10710 4320
rect 10768 4286 10784 4320
rect 10952 4286 10968 4320
rect 11026 4286 11042 4320
rect 11210 4286 11226 4320
rect 11284 4286 11300 4320
rect 11468 4286 11484 4320
rect 11542 4286 11558 4320
rect 11726 4286 11742 4320
rect 11800 4286 11816 4320
rect 11984 4286 12000 4320
rect 12058 4286 12074 4320
rect 12242 4286 12258 4320
rect 5932 4236 5966 4252
rect 5932 4044 5966 4060
rect 6190 4236 6224 4252
rect 6190 4044 6224 4060
rect 6448 4236 6482 4252
rect 6448 4044 6482 4060
rect 6706 4236 6740 4252
rect 6706 4044 6740 4060
rect 6852 4236 6886 4252
rect 6852 4044 6886 4060
rect 7110 4236 7144 4252
rect 7110 4044 7144 4060
rect 7368 4236 7402 4252
rect 7368 4044 7402 4060
rect 7626 4236 7660 4252
rect 7626 4044 7660 4060
rect 7884 4236 7918 4252
rect 7884 4044 7918 4060
rect 8142 4236 8176 4252
rect 8142 4044 8176 4060
rect 8400 4236 8434 4252
rect 8400 4044 8434 4060
rect 8658 4236 8692 4252
rect 8658 4044 8692 4060
rect 8916 4236 8950 4252
rect 8916 4044 8950 4060
rect 9174 4236 9208 4252
rect 9174 4044 9208 4060
rect 9432 4236 9466 4252
rect 9432 4044 9466 4060
rect 9690 4236 9724 4252
rect 9690 4044 9724 4060
rect 9948 4236 9982 4252
rect 9948 4044 9982 4060
rect 10206 4236 10240 4252
rect 10206 4044 10240 4060
rect 10464 4236 10498 4252
rect 10464 4044 10498 4060
rect 10722 4236 10756 4252
rect 10722 4044 10756 4060
rect 10980 4236 11014 4252
rect 10980 4044 11014 4060
rect 11238 4236 11272 4252
rect 11238 4044 11272 4060
rect 11496 4236 11530 4252
rect 11496 4044 11530 4060
rect 11754 4236 11788 4252
rect 11754 4044 11788 4060
rect 12012 4236 12046 4252
rect 12012 4044 12046 4060
rect 12270 4236 12304 4252
rect 12270 4044 12304 4060
rect 5978 3976 5994 4010
rect 6162 3976 6178 4010
rect 6236 3976 6252 4010
rect 6420 3976 6436 4010
rect 6494 3976 6510 4010
rect 6678 3976 6694 4010
rect 6898 3976 6914 4010
rect 7082 3976 7098 4010
rect 7156 3976 7172 4010
rect 7340 3976 7356 4010
rect 7414 3976 7430 4010
rect 7598 3976 7614 4010
rect 7672 3976 7688 4010
rect 7856 3976 7872 4010
rect 7930 3976 7946 4010
rect 8114 3976 8130 4010
rect 8188 3976 8204 4010
rect 8372 3976 8388 4010
rect 8446 3976 8462 4010
rect 8630 3976 8646 4010
rect 8704 3976 8720 4010
rect 8888 3976 8904 4010
rect 8962 3976 8978 4010
rect 9146 3976 9162 4010
rect 9220 3976 9236 4010
rect 9404 3976 9420 4010
rect 9478 3976 9494 4010
rect 9662 3976 9678 4010
rect 9736 3976 9752 4010
rect 9920 3976 9936 4010
rect 9994 3976 10010 4010
rect 10178 3976 10194 4010
rect 10252 3976 10268 4010
rect 10436 3976 10452 4010
rect 10510 3976 10526 4010
rect 10694 3976 10710 4010
rect 10768 3976 10784 4010
rect 10952 3976 10968 4010
rect 11026 3976 11042 4010
rect 11210 3976 11226 4010
rect 11284 3976 11300 4010
rect 11468 3976 11484 4010
rect 11542 3976 11558 4010
rect 11726 3976 11742 4010
rect 11800 3976 11816 4010
rect 11984 3976 12000 4010
rect 12058 3976 12074 4010
rect 12242 3976 12258 4010
rect 5816 3910 5850 3972
rect 12502 3910 12536 3972
rect 5816 3876 5912 3910
rect 12440 3876 12536 3910
rect 4163 3697 4197 3723
rect 243 3663 303 3697
rect 4137 3663 4197 3697
rect 17050 3562 17146 3596
rect 17304 3562 17400 3596
rect 17050 3500 17084 3562
rect 203 3303 263 3337
rect 3297 3303 3357 3337
rect 203 3277 237 3303
rect 3323 3277 3357 3303
rect 414 3107 430 3141
rect 598 3107 614 3141
rect 794 3107 810 3141
rect 978 3107 994 3141
rect 1052 3107 1068 3141
rect 1236 3107 1252 3141
rect 1310 3107 1326 3141
rect 1494 3107 1510 3141
rect 1568 3107 1584 3141
rect 1752 3107 1768 3141
rect 1826 3107 1842 3141
rect 2010 3107 2026 3141
rect 2084 3107 2100 3141
rect 2268 3107 2284 3141
rect 2342 3107 2358 3141
rect 2526 3107 2542 3141
rect 2600 3107 2616 3141
rect 2784 3107 2800 3141
rect 2974 3107 2990 3141
rect 3158 3107 3174 3141
rect 368 3048 402 3064
rect 368 2656 402 2672
rect 626 3048 660 3064
rect 626 2656 660 2672
rect 748 3048 782 3064
rect 748 2656 782 2672
rect 1006 3048 1040 3064
rect 1006 2656 1040 2672
rect 1264 3048 1298 3064
rect 1264 2656 1298 2672
rect 1522 3048 1556 3064
rect 1522 2656 1556 2672
rect 1780 3048 1814 3064
rect 1780 2656 1814 2672
rect 2038 3048 2072 3064
rect 2038 2656 2072 2672
rect 2296 3048 2330 3064
rect 2296 2656 2330 2672
rect 2554 3048 2588 3064
rect 2554 2656 2588 2672
rect 2812 3048 2846 3064
rect 2812 2656 2846 2672
rect 2928 3048 2962 3064
rect 2928 2656 2962 2672
rect 3186 3048 3220 3064
rect 14598 2995 14627 3029
rect 14661 2995 14719 3029
rect 14753 2995 14811 3029
rect 14845 2995 14903 3029
rect 14937 2995 14995 3029
rect 15029 2995 15087 3029
rect 15121 2995 15179 3029
rect 15213 2995 15271 3029
rect 15305 2995 15363 3029
rect 15397 2995 15455 3029
rect 15489 2995 15547 3029
rect 15581 2995 15639 3029
rect 15673 2995 15731 3029
rect 15765 2995 15823 3029
rect 15857 2995 15915 3029
rect 15949 2995 16007 3029
rect 16041 2995 16099 3029
rect 16133 2995 16191 3029
rect 16225 2995 16283 3029
rect 16317 2995 16375 3029
rect 16409 2995 16467 3029
rect 16501 2995 16559 3029
rect 16593 2995 16651 3029
rect 16685 2995 16714 3029
rect 14420 2960 14520 2970
rect 3186 2656 3220 2672
rect 414 2579 430 2613
rect 598 2579 614 2613
rect 794 2579 810 2613
rect 978 2579 994 2613
rect 1052 2579 1068 2613
rect 1236 2579 1252 2613
rect 1310 2579 1326 2613
rect 1494 2579 1510 2613
rect 1568 2579 1584 2613
rect 1752 2579 1768 2613
rect 1826 2579 1842 2613
rect 2010 2579 2026 2613
rect 2084 2579 2100 2613
rect 2268 2579 2284 2613
rect 2342 2579 2358 2613
rect 2526 2579 2542 2613
rect 2600 2579 2616 2613
rect 2784 2579 2800 2613
rect 2974 2579 2990 2613
rect 3158 2579 3174 2613
rect 203 2377 237 2403
rect 14420 2910 14430 2960
rect 14500 2910 14520 2960
rect 14420 2880 14520 2910
rect 14616 2945 14667 2961
rect 14616 2911 14633 2945
rect 14616 2877 14667 2911
rect 14701 2929 14767 2995
rect 14701 2895 14717 2929
rect 14751 2895 14767 2929
rect 14801 2945 14835 2961
rect 14616 2843 14633 2877
rect 14801 2877 14835 2911
rect 14667 2843 14766 2861
rect 14616 2827 14766 2843
rect 14616 2740 14686 2793
rect 14616 2680 14620 2740
rect 14660 2717 14686 2740
rect 14664 2683 14686 2717
rect 14660 2680 14686 2683
rect 14616 2663 14686 2680
rect 14720 2732 14766 2827
rect 14720 2723 14732 2732
rect 14754 2689 14766 2698
rect 14720 2629 14766 2689
rect 14616 2595 14766 2629
rect 14616 2587 14667 2595
rect 14616 2553 14633 2587
rect 14801 2587 14835 2825
rect 14869 2801 14934 2958
rect 14968 2953 15018 2995
rect 14968 2919 14984 2953
rect 14968 2903 15018 2919
rect 15052 2945 15102 2961
rect 15052 2911 15068 2945
rect 15052 2895 15102 2911
rect 15145 2951 15281 2961
rect 15145 2917 15161 2951
rect 15195 2917 15281 2951
rect 15396 2943 15462 2995
rect 15589 2953 15663 2995
rect 15145 2895 15281 2917
rect 15052 2869 15086 2895
rect 15007 2835 15086 2869
rect 15120 2859 15213 2861
rect 14881 2778 14973 2801
rect 14881 2744 14939 2778
rect 14881 2650 14973 2744
rect 14881 2610 14900 2650
rect 14960 2610 14973 2650
rect 14881 2591 14973 2610
rect 14616 2537 14667 2553
rect 14701 2527 14717 2561
rect 14751 2527 14767 2561
rect 15007 2563 15041 2835
rect 15120 2833 15179 2859
rect 15154 2825 15179 2833
rect 15154 2799 15213 2825
rect 15120 2783 15213 2799
rect 15075 2723 15145 2745
rect 15075 2689 15087 2723
rect 15121 2689 15145 2723
rect 15075 2671 15145 2689
rect 15075 2637 15098 2671
rect 15132 2637 15145 2671
rect 15075 2621 15145 2637
rect 15179 2665 15213 2783
rect 15247 2739 15281 2895
rect 15315 2927 15349 2943
rect 15396 2909 15412 2943
rect 15446 2909 15462 2943
rect 15496 2927 15530 2943
rect 15315 2875 15349 2893
rect 15589 2919 15609 2953
rect 15643 2919 15663 2953
rect 15589 2903 15663 2919
rect 15697 2945 15731 2961
rect 15496 2875 15530 2893
rect 15315 2841 15530 2875
rect 15697 2869 15731 2911
rect 15778 2952 15952 2961
rect 15778 2918 15794 2952
rect 15828 2918 15952 2952
rect 15778 2893 15952 2918
rect 15986 2953 16036 2995
rect 16020 2919 16036 2953
rect 16140 2953 16284 2995
rect 15986 2903 16036 2919
rect 16070 2927 16104 2943
rect 15619 2835 15731 2869
rect 15619 2807 15653 2835
rect 15353 2773 15369 2807
rect 15403 2773 15653 2807
rect 15792 2825 15803 2859
rect 15837 2833 15884 2859
rect 15792 2801 15834 2825
rect 15247 2719 15585 2739
rect 15247 2705 15551 2719
rect 15179 2631 15200 2665
rect 15234 2631 15250 2665
rect 15179 2621 15250 2631
rect 15284 2563 15318 2705
rect 15359 2655 15455 2671
rect 15393 2621 15431 2655
rect 15489 2637 15517 2671
rect 15551 2669 15585 2685
rect 15465 2621 15517 2637
rect 15619 2635 15653 2773
rect 14801 2537 14835 2553
rect 14701 2485 14767 2527
rect 14907 2523 14923 2557
rect 14957 2523 14973 2557
rect 15007 2529 15056 2563
rect 15090 2529 15106 2563
rect 15147 2529 15163 2563
rect 15197 2529 15318 2563
rect 15493 2561 15559 2577
rect 14907 2485 14973 2523
rect 15493 2527 15509 2561
rect 15543 2527 15559 2561
rect 15493 2485 15559 2527
rect 15601 2557 15653 2635
rect 15691 2799 15834 2801
rect 15868 2799 15884 2833
rect 15918 2817 15952 2893
rect 16140 2919 16156 2953
rect 16190 2919 16234 2953
rect 16268 2919 16284 2953
rect 16318 2945 16399 2961
rect 16550 2953 16584 2995
rect 16070 2885 16104 2893
rect 16352 2911 16399 2945
rect 16070 2851 16230 2885
rect 15691 2767 15826 2799
rect 15918 2783 16112 2817
rect 16146 2783 16162 2817
rect 15691 2659 15733 2767
rect 15918 2765 15952 2783
rect 15691 2625 15699 2659
rect 15691 2609 15733 2625
rect 15767 2723 15837 2733
rect 15767 2707 15803 2723
rect 15767 2673 15795 2707
rect 15829 2673 15837 2689
rect 15767 2609 15837 2673
rect 15871 2731 15952 2765
rect 15871 2575 15905 2731
rect 16019 2718 16127 2749
rect 16196 2733 16230 2851
rect 16318 2877 16399 2911
rect 16352 2843 16399 2877
rect 16318 2809 16399 2843
rect 16352 2775 16399 2809
rect 16318 2759 16399 2775
rect 16196 2727 16285 2733
rect 16053 2709 16127 2718
rect 15939 2681 15983 2697
rect 15973 2647 15983 2681
rect 16019 2675 16035 2684
rect 16069 2675 16127 2709
rect 15939 2641 15983 2647
rect 16079 2655 16127 2675
rect 15939 2607 16045 2641
rect 15715 2561 15905 2575
rect 15601 2523 15621 2557
rect 15655 2523 15671 2557
rect 15715 2527 15731 2561
rect 15765 2527 15905 2561
rect 15715 2519 15905 2527
rect 15939 2557 15977 2573
rect 15939 2523 15943 2557
rect 16011 2561 16045 2607
rect 16113 2621 16127 2655
rect 16079 2595 16127 2621
rect 16161 2717 16285 2727
rect 16161 2683 16235 2717
rect 16269 2683 16285 2717
rect 16161 2667 16285 2683
rect 16161 2632 16226 2667
rect 16333 2633 16399 2759
rect 16161 2577 16225 2632
rect 16011 2543 16161 2561
rect 16195 2543 16225 2577
rect 16011 2527 16225 2543
rect 16265 2600 16299 2622
rect 15939 2485 15977 2523
rect 16265 2485 16299 2566
rect 16333 2620 16349 2633
rect 16383 2620 16399 2633
rect 16437 2919 16453 2953
rect 16487 2919 16503 2953
rect 16437 2885 16503 2919
rect 16437 2851 16453 2885
rect 16487 2851 16503 2885
rect 16437 2733 16503 2851
rect 16550 2885 16584 2919
rect 16550 2817 16584 2851
rect 16550 2767 16584 2783
rect 16634 2917 16685 2933
rect 16668 2883 16685 2917
rect 16634 2849 16685 2883
rect 16668 2815 16685 2849
rect 16634 2757 16685 2815
rect 16437 2717 16609 2733
rect 16437 2683 16575 2717
rect 16437 2667 16609 2683
rect 16643 2720 16685 2757
rect 17366 3500 17400 3562
rect 17192 3460 17208 3494
rect 17242 3460 17258 3494
rect 17164 3401 17198 3417
rect 17164 2809 17198 2825
rect 17252 3401 17286 3417
rect 17252 2809 17286 2825
rect 17192 2732 17208 2766
rect 17242 2732 17258 2766
rect 16643 2680 16650 2720
rect 16333 2560 16340 2620
rect 16437 2587 16487 2667
rect 16643 2627 16685 2680
rect 17050 2664 17084 2726
rect 17366 2664 17400 2726
rect 17050 2630 17146 2664
rect 17304 2630 17400 2664
rect 16634 2611 16685 2627
rect 16333 2531 16349 2560
rect 16383 2531 16399 2560
rect 16437 2553 16453 2587
rect 16437 2537 16487 2553
rect 16550 2581 16584 2604
rect 16333 2523 16399 2531
rect 16550 2485 16584 2547
rect 16668 2577 16685 2611
rect 16634 2521 16685 2577
rect 14598 2451 14627 2485
rect 14661 2451 14719 2485
rect 14753 2451 14811 2485
rect 14845 2451 14903 2485
rect 14937 2451 14995 2485
rect 15029 2451 15087 2485
rect 15121 2451 15179 2485
rect 15213 2451 15271 2485
rect 15305 2451 15363 2485
rect 15397 2451 15455 2485
rect 15489 2451 15547 2485
rect 15581 2451 15639 2485
rect 15673 2451 15731 2485
rect 15765 2451 15823 2485
rect 15857 2451 15915 2485
rect 15949 2451 16007 2485
rect 16041 2451 16099 2485
rect 16133 2451 16191 2485
rect 16225 2451 16283 2485
rect 16317 2451 16375 2485
rect 16409 2451 16467 2485
rect 16501 2451 16559 2485
rect 16593 2451 16651 2485
rect 16685 2451 16714 2485
rect 17050 2474 17146 2508
rect 17304 2474 17400 2508
rect 3323 2377 3357 2403
rect 203 2343 263 2377
rect 3297 2343 3357 2377
rect 17050 2412 17084 2474
rect 17366 2412 17400 2474
rect 17192 2372 17208 2406
rect 17242 2372 17258 2406
rect 17164 2322 17198 2338
rect 17164 2130 17198 2146
rect 17252 2322 17286 2338
rect 17252 2130 17286 2146
rect 17192 2062 17208 2096
rect 17242 2062 17258 2096
rect 36 2010 132 2044
rect 3260 2010 3356 2044
rect 36 1948 70 2010
rect 3322 1948 3356 2010
rect 17050 1994 17084 2056
rect 17366 1994 17400 2056
rect 17050 1960 17146 1994
rect 17304 1960 17400 1994
rect 218 1910 234 1944
rect 402 1910 418 1944
rect 598 1910 614 1944
rect 782 1910 798 1944
rect 978 1910 994 1944
rect 1162 1910 1178 1944
rect 1358 1910 1374 1944
rect 1542 1910 1558 1944
rect 1738 1910 1754 1944
rect 1922 1910 1938 1944
rect 2118 1910 2134 1944
rect 2302 1910 2318 1944
rect 2498 1910 2514 1944
rect 2682 1910 2698 1944
rect 2878 1910 2894 1944
rect 3062 1910 3078 1944
rect 172 1860 206 1876
rect 172 1668 206 1684
rect 430 1860 464 1876
rect 430 1668 464 1684
rect 552 1860 586 1876
rect 552 1668 586 1684
rect 810 1860 844 1876
rect 810 1668 844 1684
rect 932 1860 966 1876
rect 932 1668 966 1684
rect 1190 1860 1224 1876
rect 1190 1668 1224 1684
rect 1312 1860 1346 1876
rect 1312 1668 1346 1684
rect 1570 1860 1604 1876
rect 1570 1668 1604 1684
rect 1692 1860 1726 1876
rect 1692 1668 1726 1684
rect 1950 1860 1984 1876
rect 1950 1668 1984 1684
rect 2072 1860 2106 1876
rect 2072 1668 2106 1684
rect 2330 1860 2364 1876
rect 2330 1668 2364 1684
rect 2452 1860 2486 1876
rect 2452 1668 2486 1684
rect 2710 1860 2744 1876
rect 2710 1668 2744 1684
rect 2832 1860 2866 1876
rect 2832 1668 2866 1684
rect 3090 1860 3124 1876
rect 3090 1668 3124 1684
rect 218 1600 234 1634
rect 402 1600 418 1634
rect 598 1600 614 1634
rect 782 1600 798 1634
rect 978 1600 994 1634
rect 1162 1600 1178 1634
rect 1358 1600 1374 1634
rect 1542 1600 1558 1634
rect 1738 1600 1754 1634
rect 1922 1600 1938 1634
rect 2118 1600 2134 1634
rect 2302 1600 2318 1634
rect 2498 1600 2514 1634
rect 2682 1600 2698 1634
rect 2878 1600 2894 1634
rect 3062 1600 3078 1634
rect 218 1492 234 1526
rect 402 1492 418 1526
rect 598 1492 614 1526
rect 782 1492 798 1526
rect 978 1492 994 1526
rect 1162 1492 1178 1526
rect 1358 1492 1374 1526
rect 1542 1492 1558 1526
rect 1738 1492 1754 1526
rect 1922 1492 1938 1526
rect 2118 1492 2134 1526
rect 2302 1492 2318 1526
rect 2498 1492 2514 1526
rect 2682 1492 2698 1526
rect 2878 1492 2894 1526
rect 3062 1492 3078 1526
rect 172 1442 206 1458
rect 172 1250 206 1266
rect 430 1442 464 1458
rect 430 1250 464 1266
rect 552 1442 586 1458
rect 552 1250 586 1266
rect 810 1442 844 1458
rect 810 1250 844 1266
rect 932 1442 966 1458
rect 932 1250 966 1266
rect 1190 1442 1224 1458
rect 1190 1250 1224 1266
rect 1312 1442 1346 1458
rect 1312 1250 1346 1266
rect 1570 1442 1604 1458
rect 1570 1250 1604 1266
rect 1692 1442 1726 1458
rect 1692 1250 1726 1266
rect 1950 1442 1984 1458
rect 1950 1250 1984 1266
rect 2072 1442 2106 1458
rect 2072 1250 2106 1266
rect 2330 1442 2364 1458
rect 2330 1250 2364 1266
rect 2452 1442 2486 1458
rect 2452 1250 2486 1266
rect 2710 1442 2744 1458
rect 2710 1250 2744 1266
rect 2832 1442 2866 1458
rect 2832 1250 2866 1266
rect 3090 1442 3124 1458
rect 3090 1250 3124 1266
rect 218 1182 234 1216
rect 402 1182 418 1216
rect 598 1182 614 1216
rect 782 1182 798 1216
rect 978 1182 994 1216
rect 1162 1182 1178 1216
rect 1358 1182 1374 1216
rect 1542 1182 1558 1216
rect 1738 1182 1754 1216
rect 1922 1182 1938 1216
rect 2118 1182 2134 1216
rect 2302 1182 2318 1216
rect 2498 1182 2514 1216
rect 2682 1182 2698 1216
rect 2878 1182 2894 1216
rect 3062 1182 3078 1216
rect 218 1074 234 1108
rect 402 1074 418 1108
rect 598 1074 614 1108
rect 782 1074 798 1108
rect 978 1074 994 1108
rect 1162 1074 1178 1108
rect 1358 1074 1374 1108
rect 1542 1074 1558 1108
rect 1738 1074 1754 1108
rect 1922 1074 1938 1108
rect 2118 1074 2134 1108
rect 2302 1074 2318 1108
rect 2498 1074 2514 1108
rect 2682 1074 2698 1108
rect 2878 1074 2894 1108
rect 3062 1074 3078 1108
rect 172 1024 206 1040
rect 172 832 206 848
rect 430 1024 464 1040
rect 430 832 464 848
rect 552 1024 586 1040
rect 552 832 586 848
rect 810 1024 844 1040
rect 810 832 844 848
rect 932 1024 966 1040
rect 932 832 966 848
rect 1190 1024 1224 1040
rect 1190 832 1224 848
rect 1312 1024 1346 1040
rect 1312 832 1346 848
rect 1570 1024 1604 1040
rect 1570 832 1604 848
rect 1692 1024 1726 1040
rect 1692 832 1726 848
rect 1950 1024 1984 1040
rect 1950 832 1984 848
rect 2072 1024 2106 1040
rect 2072 832 2106 848
rect 2330 1024 2364 1040
rect 2330 832 2364 848
rect 2452 1024 2486 1040
rect 2452 832 2486 848
rect 2710 1024 2744 1040
rect 2710 832 2744 848
rect 2832 1024 2866 1040
rect 2832 832 2866 848
rect 3090 1024 3124 1040
rect 3090 832 3124 848
rect 218 764 234 798
rect 402 764 418 798
rect 598 764 614 798
rect 782 764 798 798
rect 978 764 994 798
rect 1162 764 1178 798
rect 1358 764 1374 798
rect 1542 764 1558 798
rect 1738 764 1754 798
rect 1922 764 1938 798
rect 2118 764 2134 798
rect 2302 764 2318 798
rect 2498 764 2514 798
rect 2682 764 2698 798
rect 2878 764 2894 798
rect 3062 764 3078 798
rect 218 656 234 690
rect 402 656 418 690
rect 598 656 614 690
rect 782 656 798 690
rect 978 656 994 690
rect 1162 656 1178 690
rect 1358 656 1374 690
rect 1542 656 1558 690
rect 1738 656 1754 690
rect 1922 656 1938 690
rect 2118 656 2134 690
rect 2302 656 2318 690
rect 2498 656 2514 690
rect 2682 656 2698 690
rect 2878 656 2894 690
rect 3062 656 3078 690
rect 172 606 206 622
rect 172 414 206 430
rect 430 606 464 622
rect 430 414 464 430
rect 552 606 586 622
rect 552 414 586 430
rect 810 606 844 622
rect 810 414 844 430
rect 932 606 966 622
rect 932 414 966 430
rect 1190 606 1224 622
rect 1190 414 1224 430
rect 1312 606 1346 622
rect 1312 414 1346 430
rect 1570 606 1604 622
rect 1570 414 1604 430
rect 1692 606 1726 622
rect 1692 414 1726 430
rect 1950 606 1984 622
rect 1950 414 1984 430
rect 2072 606 2106 622
rect 2072 414 2106 430
rect 2330 606 2364 622
rect 2330 414 2364 430
rect 2452 606 2486 622
rect 2452 414 2486 430
rect 2710 606 2744 622
rect 2710 414 2744 430
rect 2832 606 2866 622
rect 2832 414 2866 430
rect 3090 606 3124 622
rect 3090 414 3124 430
rect 218 346 234 380
rect 402 346 418 380
rect 598 346 614 380
rect 782 346 798 380
rect 978 346 994 380
rect 1162 346 1178 380
rect 1358 346 1374 380
rect 1542 346 1558 380
rect 1738 346 1754 380
rect 1922 346 1938 380
rect 2118 346 2134 380
rect 2302 346 2318 380
rect 2498 346 2514 380
rect 2682 346 2698 380
rect 2878 346 2894 380
rect 3062 346 3078 380
rect 36 230 70 292
rect 3322 230 3356 292
rect 36 196 132 230
rect 3260 196 3356 230
<< viali >>
rect 6142 30835 6180 31232
rect 6142 29404 6180 29801
rect 874 10988 908 11022
rect 830 10562 864 10938
rect 918 10562 952 10938
rect 1032 10580 1066 10920
rect 874 10478 908 10512
rect 6300 6217 6420 6240
rect 6300 6183 6420 6217
rect 6300 6180 6420 6183
rect 5870 6047 6038 6081
rect 6128 6047 6296 6081
rect 6386 6047 6554 6081
rect 6644 6047 6812 6081
rect 6902 6047 7070 6081
rect 7160 6047 7328 6081
rect 7530 6047 7698 6081
rect 7910 6047 8078 6081
rect 8168 6047 8336 6081
rect 8426 6047 8594 6081
rect 8684 6047 8852 6081
rect 8942 6047 9110 6081
rect 9330 6047 9498 6081
rect 9588 6047 9756 6081
rect 9846 6047 10014 6081
rect 10104 6047 10272 6081
rect 10362 6047 10530 6081
rect 10750 6047 10918 6081
rect 11130 6047 11298 6081
rect 11388 6047 11556 6081
rect 11646 6047 11814 6081
rect 11904 6047 12072 6081
rect 12162 6047 12330 6081
rect 12420 6047 12588 6081
rect 5808 5812 5842 5988
rect 6066 5812 6100 5988
rect 6324 5812 6358 5988
rect 6582 5812 6616 5988
rect 6840 5812 6874 5988
rect 7098 5812 7132 5988
rect 7356 5812 7390 5988
rect 7468 5812 7502 5988
rect 7726 5812 7760 5988
rect 7848 5812 7882 5988
rect 8106 5812 8140 5988
rect 8364 5812 8398 5988
rect 8622 5812 8656 5988
rect 8880 5812 8914 5988
rect 9138 5812 9172 5988
rect 9268 5812 9302 5988
rect 9526 5812 9560 5988
rect 9784 5812 9818 5988
rect 10042 5812 10076 5988
rect 10300 5812 10334 5988
rect 10558 5812 10592 5988
rect 10688 5812 10722 5988
rect 10946 5812 10980 5988
rect 11068 5812 11102 5988
rect 11326 5812 11360 5988
rect 11584 5812 11618 5988
rect 11842 5812 11876 5988
rect 12100 5812 12134 5988
rect 12358 5812 12392 5988
rect 12616 5812 12650 5988
rect 5870 5719 6038 5753
rect 6128 5719 6296 5753
rect 6386 5719 6554 5753
rect 6644 5719 6812 5753
rect 6902 5719 7070 5753
rect 7160 5719 7328 5753
rect 7530 5719 7698 5753
rect 7910 5719 8078 5753
rect 8168 5719 8336 5753
rect 8426 5719 8594 5753
rect 8684 5719 8852 5753
rect 8942 5719 9110 5753
rect 9330 5719 9498 5753
rect 9588 5719 9756 5753
rect 9846 5719 10014 5753
rect 10104 5719 10272 5753
rect 10362 5719 10530 5753
rect 10750 5719 10918 5753
rect 11130 5719 11298 5753
rect 11388 5719 11556 5753
rect 11646 5719 11814 5753
rect 11904 5719 12072 5753
rect 12162 5719 12330 5753
rect 12420 5719 12588 5753
rect 14566 5337 14604 5734
rect 14732 5337 14770 5734
rect 14898 5337 14936 5734
rect 15064 5337 15102 5734
rect 15230 5337 15268 5734
rect 15396 5337 15434 5734
rect 15562 5337 15600 5734
rect 15728 5337 15766 5734
rect 16040 5337 16078 5734
rect 16206 5337 16244 5734
rect 16372 5337 16410 5734
rect 16538 5337 16576 5734
rect 16704 5337 16742 5734
rect 16870 5337 16908 5734
rect 17036 5337 17074 5734
rect 17202 5337 17240 5734
rect 840 5257 1000 5260
rect 1960 5257 2120 5260
rect 2740 5257 2900 5260
rect 3660 5257 3820 5260
rect 840 5223 1000 5257
rect 1960 5223 2120 5257
rect 2740 5223 2900 5257
rect 3660 5223 3820 5257
rect 840 5220 1000 5223
rect 1960 5220 2120 5223
rect 2740 5220 2900 5223
rect 3660 5220 3820 5223
rect 1830 5027 1998 5061
rect 2210 5027 2378 5061
rect 2590 5027 3558 5061
rect 3770 5027 3938 5061
rect 1768 4763 1802 4951
rect 2026 4763 2060 4951
rect 2148 4592 2182 4968
rect 2406 4592 2440 4968
rect 2528 4592 2562 4968
rect 3586 4592 3620 4968
rect 3708 4763 3742 4951
rect 3966 4763 4000 4951
rect 1830 4499 1998 4533
rect 2210 4499 2378 4533
rect 2590 4499 3558 4533
rect 3770 4499 3938 4533
rect 450 4347 618 4381
rect 830 4347 998 4381
rect 1088 4347 1256 4381
rect 1470 4347 1638 4381
rect 1728 4347 1896 4381
rect 1986 4347 2154 4381
rect 2244 4347 2412 4381
rect 2630 4347 2798 4381
rect 2888 4347 3056 4381
rect 3146 4347 3314 4381
rect 3404 4347 3572 4381
rect 3790 4347 3958 4381
rect 388 4083 422 4271
rect 646 4083 680 4271
rect 768 3929 802 4117
rect 1026 4083 1060 4271
rect 1284 3929 1318 4117
rect 1408 3929 1442 4117
rect 1666 4083 1700 4271
rect 1924 3929 1958 4117
rect 2182 4083 2216 4271
rect 2440 3929 2474 4117
rect 2568 3929 2602 4117
rect 2826 4083 2860 4271
rect 3084 3929 3118 4117
rect 3342 4083 3376 4271
rect 3600 3929 3634 4117
rect 3728 3929 3762 4117
rect 3986 3929 4020 4117
rect 450 3819 618 3853
rect 830 3819 998 3853
rect 1088 3819 1256 3853
rect 1470 3819 1638 3853
rect 1728 3819 1896 3853
rect 1986 3819 2154 3853
rect 2244 3819 2412 3853
rect 2630 3819 2798 3853
rect 2888 3819 3056 3853
rect 3146 3819 3314 3853
rect 3404 3819 3572 3853
rect 3790 3819 3958 3853
rect 6160 5154 6320 5160
rect 6940 5154 7100 5160
rect 7180 5154 7340 5160
rect 7960 5154 8120 5160
rect 8220 5154 8380 5160
rect 9000 5154 9160 5160
rect 9260 5154 9420 5160
rect 10020 5154 10180 5160
rect 10280 5154 10440 5160
rect 11060 5154 11220 5160
rect 6160 5120 6320 5154
rect 6940 5120 7100 5154
rect 7180 5120 7190 5154
rect 7190 5120 7340 5154
rect 7960 5120 7964 5154
rect 7964 5120 8120 5154
rect 8220 5120 8222 5154
rect 8222 5120 8380 5154
rect 9000 5120 9160 5154
rect 9260 5120 9420 5154
rect 10020 5120 10028 5154
rect 10028 5120 10180 5154
rect 10280 5120 10286 5154
rect 10286 5120 10440 5154
rect 11060 5120 11220 5154
rect 5838 4894 5872 5070
rect 6096 4894 6130 5070
rect 6354 4894 6388 5070
rect 6612 4894 6646 5070
rect 6870 4894 6904 5070
rect 7128 4894 7162 5070
rect 7386 4894 7420 5070
rect 7644 4894 7678 5070
rect 7902 4894 7936 5070
rect 8160 4894 8194 5070
rect 8418 4894 8452 5070
rect 8676 4894 8710 5070
rect 8934 4894 8968 5070
rect 9192 4894 9226 5070
rect 9450 4894 9484 5070
rect 9708 4894 9742 5070
rect 9966 4894 10000 5070
rect 10224 4894 10258 5070
rect 10482 4894 10516 5070
rect 10740 4894 10774 5070
rect 10998 4894 11032 5070
rect 11256 4894 11290 5070
rect 11514 4894 11548 5070
rect 5900 4810 6060 4840
rect 6420 4810 6580 4840
rect 6680 4810 6840 4840
rect 7440 4810 7448 4840
rect 7448 4810 7600 4840
rect 7700 4810 7706 4840
rect 7706 4810 7860 4840
rect 8480 4810 8640 4840
rect 8740 4810 8900 4840
rect 9520 4810 9680 4840
rect 9760 4810 9770 4840
rect 9770 4810 9920 4840
rect 10540 4810 10544 4840
rect 10544 4810 10700 4840
rect 10800 4810 10802 4840
rect 10802 4810 10960 4840
rect 11320 4810 11480 4840
rect 5900 4800 6060 4810
rect 6420 4800 6580 4810
rect 6680 4800 6840 4810
rect 7440 4800 7600 4810
rect 7700 4800 7860 4810
rect 8480 4800 8640 4810
rect 8740 4800 8900 4810
rect 9520 4800 9680 4810
rect 9760 4800 9920 4810
rect 10540 4800 10700 4810
rect 10800 4800 10960 4810
rect 11320 4800 11480 4810
rect 5994 4286 6162 4320
rect 6252 4286 6420 4320
rect 6510 4286 6678 4320
rect 6914 4286 7082 4320
rect 7172 4286 7340 4320
rect 7430 4286 7598 4320
rect 7688 4286 7856 4320
rect 7946 4286 8114 4320
rect 8204 4286 8372 4320
rect 8462 4286 8630 4320
rect 8720 4286 8888 4320
rect 8978 4286 9146 4320
rect 9236 4286 9404 4320
rect 9494 4286 9662 4320
rect 9752 4286 9920 4320
rect 10010 4286 10178 4320
rect 10268 4286 10436 4320
rect 10526 4286 10694 4320
rect 10784 4286 10952 4320
rect 11042 4286 11210 4320
rect 11300 4286 11468 4320
rect 11558 4286 11726 4320
rect 11816 4286 11984 4320
rect 12074 4286 12242 4320
rect 5932 4060 5966 4236
rect 6190 4060 6224 4236
rect 6448 4060 6482 4236
rect 6706 4060 6740 4236
rect 6852 4060 6886 4236
rect 7110 4060 7144 4236
rect 7368 4060 7402 4236
rect 7626 4060 7660 4236
rect 7884 4060 7918 4236
rect 8142 4060 8176 4236
rect 8400 4060 8434 4236
rect 8658 4060 8692 4236
rect 8916 4060 8950 4236
rect 9174 4060 9208 4236
rect 9432 4060 9466 4236
rect 9690 4060 9724 4236
rect 9948 4060 9982 4236
rect 10206 4060 10240 4236
rect 10464 4060 10498 4236
rect 10722 4060 10756 4236
rect 10980 4060 11014 4236
rect 11238 4060 11272 4236
rect 11496 4060 11530 4236
rect 11754 4060 11788 4236
rect 12012 4060 12046 4236
rect 12270 4060 12304 4236
rect 5994 3976 6162 4010
rect 6252 3976 6420 4010
rect 6510 3976 6678 4010
rect 6914 3976 7082 4010
rect 7172 3976 7340 4010
rect 7430 3976 7598 4010
rect 7688 3976 7856 4010
rect 7946 3976 8114 4010
rect 8204 3976 8372 4010
rect 8462 3976 8630 4010
rect 8720 3976 8888 4010
rect 8978 3976 9146 4010
rect 9236 3976 9404 4010
rect 9494 3976 9662 4010
rect 9752 3976 9920 4010
rect 10010 3976 10178 4010
rect 10268 3976 10436 4010
rect 10526 3976 10694 4010
rect 10784 3976 10952 4010
rect 11042 3976 11210 4010
rect 11300 3976 11468 4010
rect 11558 3976 11726 4010
rect 11816 3976 11984 4010
rect 12074 3976 12242 4010
rect 14566 4006 14604 4403
rect 14732 4006 14770 4403
rect 14898 4006 14936 4403
rect 15064 4006 15102 4403
rect 15230 4006 15268 4403
rect 15396 4006 15434 4403
rect 15562 4006 15600 4403
rect 15728 4006 15766 4403
rect 16040 4006 16078 4403
rect 16206 4006 16244 4403
rect 16372 4006 16410 4403
rect 16538 4006 16576 4403
rect 16704 4006 16742 4403
rect 16870 4006 16908 4403
rect 17036 4006 17074 4403
rect 17202 4006 17240 4403
rect 6040 3910 6380 3920
rect 6040 3876 6380 3910
rect 6040 3860 6380 3876
rect 430 3107 598 3141
rect 810 3107 978 3141
rect 1068 3107 1236 3141
rect 1326 3107 1494 3141
rect 1584 3107 1752 3141
rect 1842 3107 2010 3141
rect 2100 3107 2268 3141
rect 2358 3107 2526 3141
rect 2616 3107 2784 3141
rect 2990 3107 3158 3141
rect 368 2843 402 3031
rect 626 2843 660 3031
rect 748 2689 782 2877
rect 1006 2843 1040 3031
rect 1264 2689 1298 2877
rect 1522 2843 1556 3031
rect 1780 2689 1814 2877
rect 2038 2843 2072 3031
rect 2296 2689 2330 2877
rect 2554 2843 2588 3031
rect 2812 2689 2846 2877
rect 2928 2843 2962 3031
rect 3186 2843 3220 3031
rect 3280 2940 3323 3040
rect 3323 2940 3357 3040
rect 3357 2940 3360 3040
rect 14627 2995 14661 3029
rect 14719 2995 14753 3029
rect 14811 2995 14845 3029
rect 14903 2995 14937 3029
rect 14995 2995 15029 3029
rect 15087 2995 15121 3029
rect 15179 2995 15213 3029
rect 15271 2995 15305 3029
rect 15363 2995 15397 3029
rect 15455 2995 15489 3029
rect 15547 2995 15581 3029
rect 15639 2995 15673 3029
rect 15731 2995 15765 3029
rect 15823 2995 15857 3029
rect 15915 2995 15949 3029
rect 16007 2995 16041 3029
rect 16099 2995 16133 3029
rect 16191 2995 16225 3029
rect 16283 2995 16317 3029
rect 16375 2995 16409 3029
rect 16467 2995 16501 3029
rect 16559 2995 16593 3029
rect 16651 2995 16685 3029
rect 430 2579 598 2613
rect 810 2579 978 2613
rect 1068 2579 1236 2613
rect 1326 2579 1494 2613
rect 1584 2579 1752 2613
rect 1842 2579 2010 2613
rect 2100 2579 2268 2613
rect 2358 2579 2526 2613
rect 2616 2579 2784 2613
rect 2990 2579 3158 2613
rect 14430 2950 14500 2960
rect 14430 2910 14450 2950
rect 14450 2910 14490 2950
rect 14490 2910 14500 2950
rect 14620 2717 14660 2740
rect 14620 2683 14630 2717
rect 14630 2683 14660 2717
rect 14620 2680 14660 2683
rect 14720 2698 14732 2723
rect 14732 2698 14754 2723
rect 14720 2689 14754 2698
rect 14801 2843 14835 2859
rect 14801 2825 14835 2843
rect 14900 2610 14960 2650
rect 15179 2825 15213 2859
rect 15087 2689 15121 2723
rect 15803 2833 15837 2859
rect 15803 2825 15834 2833
rect 15834 2825 15837 2833
rect 15359 2621 15393 2655
rect 15431 2637 15455 2655
rect 15455 2637 15465 2655
rect 15431 2621 15465 2637
rect 15803 2707 15837 2723
rect 15803 2689 15829 2707
rect 15829 2689 15837 2707
rect 16019 2709 16053 2718
rect 16019 2684 16035 2709
rect 16035 2684 16053 2709
rect 16079 2621 16113 2655
rect 17208 3460 17242 3494
rect 17164 2825 17198 3401
rect 17252 2825 17286 3401
rect 17360 2840 17366 3400
rect 17366 2840 17400 3400
rect 17208 2732 17242 2766
rect 16650 2680 16690 2720
rect 16340 2599 16349 2620
rect 16349 2599 16383 2620
rect 16383 2599 16400 2620
rect 16340 2565 16400 2599
rect 16340 2560 16349 2565
rect 16349 2560 16383 2565
rect 16383 2560 16400 2565
rect 14627 2451 14661 2485
rect 14719 2451 14753 2485
rect 14811 2451 14845 2485
rect 14903 2451 14937 2485
rect 14995 2451 15029 2485
rect 15087 2451 15121 2485
rect 15179 2451 15213 2485
rect 15271 2451 15305 2485
rect 15363 2451 15397 2485
rect 15455 2451 15489 2485
rect 15547 2451 15581 2485
rect 15639 2451 15673 2485
rect 15731 2451 15765 2485
rect 15823 2451 15857 2485
rect 15915 2451 15949 2485
rect 16007 2451 16041 2485
rect 16099 2451 16133 2485
rect 16191 2451 16225 2485
rect 16283 2451 16317 2485
rect 16375 2451 16409 2485
rect 16467 2451 16501 2485
rect 16559 2451 16593 2485
rect 16651 2451 16685 2485
rect 17208 2372 17242 2406
rect 17164 2146 17198 2322
rect 17252 2146 17286 2322
rect 17360 2140 17366 2300
rect 17366 2140 17400 2300
rect 17208 2062 17242 2096
rect 234 1910 402 1944
rect 614 1910 782 1944
rect 994 1910 1162 1944
rect 1374 1910 1542 1944
rect 1754 1910 1922 1944
rect 2134 1910 2302 1944
rect 2514 1910 2682 1944
rect 2894 1910 3062 1944
rect 172 1684 206 1860
rect 430 1684 464 1860
rect 552 1684 586 1860
rect 810 1684 844 1860
rect 932 1684 966 1860
rect 1190 1684 1224 1860
rect 1312 1684 1346 1860
rect 1570 1684 1604 1860
rect 1692 1684 1726 1860
rect 1950 1684 1984 1860
rect 2072 1684 2106 1860
rect 2330 1684 2364 1860
rect 2452 1684 2486 1860
rect 2710 1684 2744 1860
rect 2832 1684 2866 1860
rect 3090 1684 3124 1860
rect 234 1600 402 1634
rect 614 1600 782 1634
rect 994 1600 1162 1634
rect 1374 1600 1542 1634
rect 1754 1600 1922 1634
rect 2134 1600 2302 1634
rect 2514 1600 2682 1634
rect 2894 1600 3062 1634
rect 234 1492 402 1526
rect 614 1492 782 1526
rect 994 1492 1162 1526
rect 1374 1492 1542 1526
rect 1754 1492 1922 1526
rect 2134 1492 2302 1526
rect 2514 1492 2682 1526
rect 2894 1492 3062 1526
rect 172 1266 206 1442
rect 430 1266 464 1442
rect 552 1266 586 1442
rect 810 1266 844 1442
rect 932 1266 966 1442
rect 1190 1266 1224 1442
rect 1312 1266 1346 1442
rect 1570 1266 1604 1442
rect 1692 1266 1726 1442
rect 1950 1266 1984 1442
rect 2072 1266 2106 1442
rect 2330 1266 2364 1442
rect 2452 1266 2486 1442
rect 2710 1266 2744 1442
rect 2832 1266 2866 1442
rect 3090 1266 3124 1442
rect 234 1182 402 1216
rect 614 1182 782 1216
rect 994 1182 1162 1216
rect 1374 1182 1542 1216
rect 1754 1182 1922 1216
rect 2134 1182 2302 1216
rect 2514 1182 2682 1216
rect 2894 1182 3062 1216
rect 234 1074 402 1108
rect 614 1074 782 1108
rect 994 1074 1162 1108
rect 1374 1074 1542 1108
rect 1754 1074 1922 1108
rect 2134 1074 2302 1108
rect 2514 1074 2682 1108
rect 2894 1074 3062 1108
rect 172 848 206 1024
rect 430 848 464 1024
rect 552 848 586 1024
rect 810 848 844 1024
rect 932 848 966 1024
rect 1190 848 1224 1024
rect 1312 848 1346 1024
rect 1570 848 1604 1024
rect 1692 848 1726 1024
rect 1950 848 1984 1024
rect 2072 848 2106 1024
rect 2330 848 2364 1024
rect 2452 848 2486 1024
rect 2710 848 2744 1024
rect 2832 848 2866 1024
rect 3090 848 3124 1024
rect 234 764 402 798
rect 614 764 782 798
rect 994 764 1162 798
rect 1374 764 1542 798
rect 1754 764 1922 798
rect 2134 764 2302 798
rect 2514 764 2682 798
rect 2894 764 3062 798
rect 234 656 402 690
rect 614 656 782 690
rect 994 656 1162 690
rect 1374 656 1542 690
rect 1754 656 1922 690
rect 2134 656 2302 690
rect 2514 656 2682 690
rect 2894 656 3062 690
rect 172 430 206 606
rect 430 430 464 606
rect 552 430 586 606
rect 810 430 844 606
rect 932 430 966 606
rect 1190 430 1224 606
rect 1312 430 1346 606
rect 1570 430 1604 606
rect 1692 430 1726 606
rect 1950 430 1984 606
rect 2072 430 2106 606
rect 2330 430 2364 606
rect 2452 430 2486 606
rect 2710 430 2744 606
rect 2832 430 2866 606
rect 3090 430 3124 606
rect 234 346 402 380
rect 614 346 782 380
rect 994 346 1162 380
rect 1374 346 1542 380
rect 1754 346 1922 380
rect 2134 346 2302 380
rect 2514 346 2682 380
rect 2894 346 3062 380
rect 220 230 440 240
rect 1100 230 1320 240
rect 2020 230 2240 240
rect 2860 230 3080 240
rect 220 200 440 230
rect 1100 200 1320 230
rect 2020 200 2240 230
rect 2860 200 3080 230
<< metal1 >>
rect 6000 33780 7320 33820
rect 6000 33500 6940 33780
rect 7260 33500 7320 33780
rect 6000 33480 7320 33500
rect 6040 33160 6240 33480
rect 6040 33060 6260 33160
rect 5850 32440 5860 33060
rect 6460 32440 6470 33060
rect 5830 30800 5840 31400
rect 6440 30800 6450 31400
rect 6136 29801 6186 29813
rect 6136 29404 6142 29801
rect 6180 29404 6186 29801
rect 6136 29392 6186 29404
rect -80 11320 1580 11460
rect 1760 11320 1780 11460
rect -80 11300 1780 11320
rect -80 11260 120 11300
rect 860 11022 920 11300
rect 860 10988 874 11022
rect 908 10988 920 11022
rect 860 10980 920 10988
rect 210 10920 220 10980
rect -320 10720 220 10920
rect 210 10660 220 10720
rect 500 10920 510 10980
rect 824 10938 870 10950
rect 824 10920 830 10938
rect 500 10720 830 10920
rect 500 10660 510 10720
rect 824 10562 830 10720
rect 864 10562 870 10938
rect 824 10550 870 10562
rect 912 10938 958 10950
rect 912 10562 918 10938
rect 952 10920 958 10938
rect 1026 10920 1072 10932
rect 952 10580 1032 10920
rect 1066 10580 1240 10920
rect 952 10562 958 10580
rect 1026 10568 1240 10580
rect 912 10550 958 10562
rect 860 10512 920 10520
rect 860 10478 874 10512
rect 908 10478 920 10512
rect 860 10460 920 10478
rect 1040 6560 1240 10568
rect 1550 6760 13100 6780
rect 1550 6560 1560 6760
rect 1760 6560 12880 6760
rect 13080 6560 13100 6760
rect 1030 6400 1040 6560
rect 1220 6400 1240 6560
rect 1040 6380 1240 6400
rect 6280 6420 6480 6440
rect 6280 6280 6300 6420
rect 6460 6280 6480 6420
rect 6280 6260 6480 6280
rect 6050 6180 6060 6260
rect 6120 6240 6580 6260
rect 6120 6200 6300 6240
rect 6120 6180 6130 6200
rect 6288 6180 6300 6200
rect 6420 6200 6580 6240
rect 6420 6180 6432 6200
rect 6570 6180 6580 6200
rect 6640 6180 7080 6260
rect 7140 6200 7460 6260
rect 7520 6200 8100 6260
rect 7140 6180 8100 6200
rect 8160 6180 8620 6260
rect 8680 6180 9120 6260
rect 9180 6180 9520 6260
rect 9580 6180 10020 6260
rect 10080 6180 10540 6260
rect 10600 6180 10680 6260
rect 10740 6180 11320 6260
rect 11380 6180 11840 6260
rect 11900 6180 12360 6260
rect 12420 6180 12430 6260
rect 6288 6174 6432 6180
rect 5858 6081 6050 6087
rect 5858 6080 5870 6081
rect 5840 6047 5870 6080
rect 6038 6080 6050 6081
rect 6116 6081 6308 6087
rect 6038 6047 6060 6080
rect 5840 6000 6060 6047
rect 6116 6047 6128 6081
rect 6296 6047 6308 6081
rect 6116 6041 6308 6047
rect 6374 6081 6566 6087
rect 6374 6047 6386 6081
rect 6554 6047 6566 6081
rect 6374 6041 6566 6047
rect 6632 6081 6824 6087
rect 6632 6047 6644 6081
rect 6812 6047 6824 6081
rect 6632 6041 6824 6047
rect 6890 6081 7082 6087
rect 6890 6047 6902 6081
rect 7070 6047 7082 6081
rect 6890 6041 7082 6047
rect 7148 6081 7340 6087
rect 7148 6047 7160 6081
rect 7328 6047 7340 6081
rect 7148 6041 7340 6047
rect 7518 6081 7710 6087
rect 7518 6047 7530 6081
rect 7698 6047 7710 6081
rect 7518 6041 7710 6047
rect 7898 6081 8090 6087
rect 7898 6047 7910 6081
rect 8078 6047 8090 6081
rect 7898 6041 8090 6047
rect 8156 6081 8348 6087
rect 8156 6047 8168 6081
rect 8336 6047 8348 6081
rect 8156 6041 8348 6047
rect 8414 6081 8606 6087
rect 8414 6047 8426 6081
rect 8594 6047 8606 6081
rect 8414 6041 8606 6047
rect 8672 6081 8864 6087
rect 8672 6047 8684 6081
rect 8852 6047 8864 6081
rect 8672 6041 8864 6047
rect 8930 6081 9122 6087
rect 8930 6047 8942 6081
rect 9110 6047 9122 6081
rect 8930 6041 9122 6047
rect 9318 6081 9510 6087
rect 9318 6047 9330 6081
rect 9498 6047 9510 6081
rect 9318 6041 9510 6047
rect 9576 6081 9768 6087
rect 9576 6047 9588 6081
rect 9756 6047 9768 6081
rect 9576 6041 9768 6047
rect 9834 6081 10026 6087
rect 9834 6047 9846 6081
rect 10014 6047 10026 6081
rect 9834 6041 10026 6047
rect 10092 6081 10284 6087
rect 10092 6047 10104 6081
rect 10272 6047 10284 6081
rect 10092 6041 10284 6047
rect 10350 6081 10542 6087
rect 10350 6047 10362 6081
rect 10530 6047 10542 6081
rect 10350 6041 10542 6047
rect 10738 6081 10930 6087
rect 10738 6047 10750 6081
rect 10918 6047 10930 6081
rect 10738 6041 10930 6047
rect 11118 6081 11310 6087
rect 11118 6047 11130 6081
rect 11298 6047 11310 6081
rect 11118 6041 11310 6047
rect 11376 6081 11568 6087
rect 11376 6047 11388 6081
rect 11556 6047 11568 6081
rect 11376 6041 11568 6047
rect 11634 6081 11826 6087
rect 11634 6047 11646 6081
rect 11814 6047 11826 6081
rect 11634 6041 11826 6047
rect 11892 6081 12084 6087
rect 11892 6047 11904 6081
rect 12072 6047 12084 6081
rect 11892 6041 12084 6047
rect 12150 6081 12342 6087
rect 12150 6047 12162 6081
rect 12330 6047 12342 6081
rect 12408 6081 12600 6087
rect 12408 6080 12420 6081
rect 12150 6041 12342 6047
rect 12400 6047 12420 6080
rect 12588 6080 12600 6081
rect 12588 6047 12620 6080
rect 12400 6000 12620 6047
rect 5800 5988 6060 6000
rect 5800 5820 5808 5988
rect 5802 5812 5808 5820
rect 5842 5812 6060 5988
rect 5802 5800 6060 5812
rect 6120 5800 6130 6000
rect 6290 5800 6300 6000
rect 6360 5800 6370 6000
rect 6570 5800 6580 6000
rect 6640 5800 6650 6000
rect 6810 5800 6820 6000
rect 6880 5800 6890 6000
rect 7070 5800 7080 6000
rect 7140 5800 7150 6000
rect 7330 5800 7340 6000
rect 7400 5800 7410 6000
rect 7450 5800 7460 6000
rect 7520 5800 7530 6000
rect 7690 5800 7700 6000
rect 7760 5800 7770 6000
rect 7830 5800 7840 6000
rect 7900 5800 7910 6000
rect 8090 5800 8100 6000
rect 8160 5800 8170 6000
rect 8350 5800 8360 6000
rect 8420 5800 8430 6000
rect 8590 5800 8600 6000
rect 8660 5800 8670 6000
rect 8850 5800 8860 6000
rect 8920 5800 8930 6000
rect 9110 5800 9120 6000
rect 9180 5800 9190 6000
rect 9250 5800 9260 6000
rect 9320 5800 9330 6000
rect 9510 5800 9520 6000
rect 9580 5800 9590 6000
rect 9770 5800 9780 6000
rect 9840 5800 9850 6000
rect 10010 5800 10020 6000
rect 10080 5800 10090 6000
rect 10270 5800 10280 6000
rect 10340 5800 10350 6000
rect 10530 5800 10540 6000
rect 10600 5800 10610 6000
rect 10670 5800 10680 6000
rect 10740 5800 10750 6000
rect 10930 5988 11010 6000
rect 10930 5812 10946 5988
rect 10980 5812 11010 5988
rect 10930 5800 11010 5812
rect 11050 5800 11060 6000
rect 11120 5800 11130 6000
rect 11310 5800 11320 6000
rect 11380 5800 11390 6000
rect 11550 5800 11560 6000
rect 11620 5800 11630 6000
rect 11830 5800 11840 6000
rect 11900 5800 11910 6000
rect 12090 5800 12100 6000
rect 12160 5800 12170 6000
rect 12350 5988 12360 6000
rect 12420 5988 12660 6000
rect 12350 5812 12358 5988
rect 12420 5812 12616 5988
rect 12650 5812 12660 5988
rect 12350 5800 12360 5812
rect 12420 5800 12660 5812
rect 5840 5753 6060 5800
rect 7720 5760 7760 5800
rect 10790 5760 10870 5800
rect 10940 5760 11000 5800
rect 6120 5759 9120 5760
rect 9320 5759 12340 5760
rect 5840 5720 5870 5753
rect 5858 5719 5870 5720
rect 6038 5720 6060 5753
rect 6116 5753 9122 5759
rect 6038 5719 6050 5720
rect 5858 5713 6050 5719
rect 6116 5719 6128 5753
rect 6296 5720 6386 5753
rect 6296 5719 6308 5720
rect 6116 5713 6308 5719
rect 6374 5719 6386 5720
rect 6554 5720 6644 5753
rect 6554 5719 6566 5720
rect 6374 5713 6566 5719
rect 6632 5719 6644 5720
rect 6812 5720 6902 5753
rect 6812 5719 6824 5720
rect 6632 5713 6824 5719
rect 6890 5719 6902 5720
rect 7070 5720 7160 5753
rect 7070 5719 7082 5720
rect 6890 5713 7082 5719
rect 7148 5719 7160 5720
rect 7328 5720 7530 5753
rect 7328 5719 7340 5720
rect 7148 5713 7340 5719
rect 7518 5719 7530 5720
rect 7698 5720 7910 5753
rect 7698 5719 7710 5720
rect 7518 5713 7710 5719
rect 7898 5719 7910 5720
rect 8078 5720 8168 5753
rect 8078 5719 8090 5720
rect 7898 5713 8090 5719
rect 8156 5719 8168 5720
rect 8336 5720 8426 5753
rect 8336 5719 8348 5720
rect 8156 5713 8348 5719
rect 8414 5719 8426 5720
rect 8594 5720 8684 5753
rect 8594 5719 8606 5720
rect 8414 5713 8606 5719
rect 8672 5719 8684 5720
rect 8852 5720 8942 5753
rect 8852 5719 8864 5720
rect 8672 5713 8864 5719
rect 8930 5719 8942 5720
rect 9110 5719 9122 5753
rect 8930 5713 9122 5719
rect 9318 5753 12342 5759
rect 9318 5719 9330 5753
rect 9498 5720 9588 5753
rect 9498 5719 9510 5720
rect 9318 5713 9510 5719
rect 9576 5719 9588 5720
rect 9756 5720 9846 5753
rect 9756 5719 9768 5720
rect 9576 5713 9768 5719
rect 9834 5719 9846 5720
rect 10014 5720 10104 5753
rect 10014 5719 10026 5720
rect 9834 5713 10026 5719
rect 10092 5719 10104 5720
rect 10272 5720 10362 5753
rect 10272 5719 10284 5720
rect 10092 5713 10284 5719
rect 10350 5719 10362 5720
rect 10530 5740 10750 5753
rect 10530 5720 10720 5740
rect 10530 5719 10542 5720
rect 10350 5713 10542 5719
rect 10710 5680 10720 5720
rect 10918 5720 11130 5753
rect 10918 5719 10930 5720
rect 10780 5713 10930 5719
rect 11118 5719 11130 5720
rect 11298 5720 11388 5753
rect 11298 5719 11310 5720
rect 11118 5713 11310 5719
rect 11376 5719 11388 5720
rect 11556 5720 11646 5753
rect 11556 5719 11568 5720
rect 11376 5713 11568 5719
rect 11634 5719 11646 5720
rect 11814 5720 11904 5753
rect 11814 5719 11826 5720
rect 11634 5713 11826 5719
rect 11892 5719 11904 5720
rect 12072 5720 12162 5753
rect 12072 5719 12084 5720
rect 11892 5713 12084 5719
rect 12150 5719 12162 5720
rect 12330 5719 12342 5753
rect 12400 5753 12620 5800
rect 12400 5720 12420 5753
rect 12150 5713 12342 5719
rect 12408 5719 12420 5720
rect 12588 5720 12620 5753
rect 14560 5740 14610 5746
rect 14726 5740 14776 5746
rect 14540 5734 14776 5740
rect 12588 5719 12600 5720
rect 12408 5713 12600 5719
rect 10780 5680 10790 5713
rect 6280 5540 6300 5620
rect 6360 5600 6380 5620
rect 6810 5600 6820 5620
rect 6360 5540 6820 5600
rect 6880 5600 6890 5620
rect 7330 5600 7340 5620
rect 6880 5540 7220 5600
rect 7280 5540 7340 5600
rect 7400 5600 7410 5620
rect 7830 5600 7840 5620
rect 7400 5540 7840 5600
rect 7900 5600 7910 5620
rect 8350 5600 8360 5620
rect 7900 5540 8360 5600
rect 8420 5600 8430 5620
rect 8850 5600 8860 5620
rect 8420 5540 8860 5600
rect 8920 5540 8930 5620
rect 9230 5540 9240 5620
rect 9300 5600 9310 5620
rect 9750 5600 9760 5620
rect 9300 5540 9760 5600
rect 9820 5600 9830 5620
rect 10270 5600 10280 5620
rect 9820 5540 10280 5600
rect 10340 5600 10350 5620
rect 11050 5600 11060 5620
rect 10340 5540 10600 5600
rect 10660 5540 11060 5600
rect 11120 5600 11130 5620
rect 11550 5600 11560 5620
rect 11120 5540 11560 5600
rect 11620 5600 11630 5620
rect 12090 5600 12100 5620
rect 11620 5540 12100 5600
rect 12160 5540 12170 5620
rect 4360 5520 5840 5540
rect 320 5480 4240 5500
rect 320 5400 3500 5480
rect 310 5300 320 5400
rect 400 5300 1600 5400
rect 1720 5320 3500 5400
rect 4000 5400 4240 5480
rect 4000 5320 4040 5400
rect 1720 5300 4040 5320
rect 4140 5300 4240 5400
rect 4360 5340 4380 5520
rect 4560 5480 5840 5520
rect 4560 5420 6180 5480
rect 6240 5420 6250 5480
rect 4560 5340 5840 5420
rect 12600 5400 14480 5420
rect 6330 5320 6340 5380
rect 6400 5320 6700 5380
rect 6760 5320 6860 5380
rect 6920 5320 7360 5380
rect 7420 5320 7880 5380
rect 7940 5320 8400 5380
rect 8460 5320 8920 5380
rect 8980 5320 9420 5380
rect 9480 5320 9940 5380
rect 10000 5320 10460 5380
rect 10520 5320 10980 5380
rect 11040 5320 11050 5380
rect 11110 5340 11120 5400
rect 11180 5340 11600 5400
rect 11120 5320 11600 5340
rect 11660 5320 14300 5400
rect 840 5266 1000 5300
rect 1960 5266 2120 5300
rect 2740 5266 2900 5300
rect 3660 5266 3820 5300
rect 828 5260 1012 5266
rect 828 5220 840 5260
rect 1000 5220 1012 5260
rect 828 5214 1012 5220
rect 1948 5260 2132 5266
rect 1948 5220 1960 5260
rect 2120 5220 2132 5260
rect 1948 5214 2132 5220
rect 2728 5260 2912 5266
rect 2728 5220 2740 5260
rect 2900 5220 2912 5260
rect 2728 5214 2912 5220
rect 3648 5260 3832 5266
rect 3648 5220 3660 5260
rect 3820 5220 3832 5260
rect 3648 5214 3832 5220
rect 6050 5200 6060 5260
rect 6120 5200 7100 5260
rect 7160 5200 7700 5260
rect 7760 5200 8140 5260
rect 8200 5200 9160 5260
rect 9220 5200 10200 5260
rect 10260 5200 11240 5260
rect 11300 5200 11320 5260
rect 12600 5240 14300 5320
rect 14440 5240 14480 5400
rect 14540 5340 14566 5734
rect 14560 5337 14566 5340
rect 14604 5340 14732 5734
rect 14604 5337 14610 5340
rect 14560 5325 14610 5337
rect 14726 5337 14732 5340
rect 14770 5337 14776 5734
rect 14726 5325 14776 5337
rect 14892 5740 14942 5746
rect 15058 5740 15108 5746
rect 15224 5740 15274 5746
rect 15390 5740 15440 5746
rect 14892 5734 15120 5740
rect 14892 5337 14898 5734
rect 14936 5340 15064 5734
rect 14936 5337 14942 5340
rect 14892 5325 14942 5337
rect 15058 5337 15064 5340
rect 15102 5340 15120 5734
rect 15220 5734 15440 5740
rect 15220 5340 15230 5734
rect 15102 5337 15108 5340
rect 15058 5325 15108 5337
rect 15224 5337 15230 5340
rect 15268 5340 15396 5734
rect 15268 5337 15274 5340
rect 15224 5325 15274 5337
rect 15390 5337 15396 5340
rect 15434 5337 15440 5734
rect 15390 5325 15440 5337
rect 15556 5740 15606 5746
rect 15722 5740 15772 5746
rect 16034 5740 16084 5746
rect 16200 5740 16250 5746
rect 16366 5740 16416 5746
rect 16532 5740 16582 5746
rect 16698 5740 16748 5746
rect 16864 5740 16914 5746
rect 17030 5740 17080 5746
rect 17196 5740 17246 5746
rect 15556 5734 15780 5740
rect 15556 5337 15562 5734
rect 15600 5340 15728 5734
rect 15600 5337 15606 5340
rect 15556 5325 15606 5337
rect 15722 5337 15728 5340
rect 15766 5340 15780 5734
rect 16034 5734 16260 5740
rect 15766 5337 15772 5340
rect 15722 5325 15772 5337
rect 16034 5337 16040 5734
rect 16078 5340 16206 5734
rect 16078 5337 16084 5340
rect 16034 5325 16084 5337
rect 16200 5337 16206 5340
rect 16244 5340 16260 5734
rect 16366 5734 16600 5740
rect 16244 5337 16250 5340
rect 16200 5325 16250 5337
rect 16366 5337 16372 5734
rect 16410 5340 16538 5734
rect 16410 5337 16416 5340
rect 16366 5325 16416 5337
rect 16532 5337 16538 5340
rect 16576 5340 16600 5734
rect 16698 5734 16920 5740
rect 16576 5337 16582 5340
rect 16532 5325 16582 5337
rect 16698 5337 16704 5734
rect 16742 5340 16870 5734
rect 16742 5337 16748 5340
rect 16698 5325 16748 5337
rect 16864 5337 16870 5340
rect 16908 5340 16920 5734
rect 17030 5734 17260 5740
rect 16908 5337 16914 5340
rect 16864 5325 16914 5337
rect 17030 5337 17036 5734
rect 17074 5340 17202 5734
rect 17074 5337 17080 5340
rect 17030 5325 17080 5337
rect 17196 5337 17202 5340
rect 17240 5340 17260 5734
rect 17310 5700 17320 5880
rect 17500 5700 17540 5880
rect 17340 5680 17540 5700
rect 17340 5520 17460 5680
rect 17340 5440 17360 5520
rect 17460 5440 17470 5520
rect 17240 5337 17246 5340
rect 17196 5325 17246 5337
rect 12600 5220 14480 5240
rect 6148 5160 6332 5166
rect 6928 5160 7112 5166
rect 7168 5160 7352 5166
rect 7948 5160 8132 5166
rect 8208 5160 8392 5166
rect 8988 5160 9172 5166
rect 9248 5160 9432 5166
rect 10008 5160 10192 5166
rect 10268 5160 10452 5166
rect 11048 5160 11232 5166
rect 5860 5082 6100 5160
rect 6148 5120 6160 5160
rect 6320 5120 6940 5160
rect 7100 5120 7180 5160
rect 7340 5120 7960 5160
rect 8120 5120 8220 5160
rect 8380 5120 9000 5160
rect 9160 5120 9260 5160
rect 9420 5120 10020 5160
rect 10180 5120 10280 5160
rect 10440 5120 11060 5160
rect 11220 5120 11232 5160
rect 6148 5114 6332 5120
rect 6928 5114 7112 5120
rect 7168 5114 7352 5120
rect 7948 5114 8132 5120
rect 8208 5114 8392 5120
rect 8988 5114 9172 5120
rect 9248 5114 9432 5120
rect 10008 5114 10192 5120
rect 10268 5114 10452 5120
rect 11048 5114 11120 5120
rect 11110 5100 11120 5114
rect 11180 5114 11232 5120
rect 11180 5100 11190 5114
rect 11280 5082 11520 5160
rect 5832 5080 6136 5082
rect 6348 5080 6394 5082
rect 6606 5080 6652 5082
rect 6864 5080 6910 5082
rect 7122 5080 7168 5082
rect 7380 5080 7426 5082
rect 7638 5080 7684 5082
rect 7896 5080 7942 5082
rect 8154 5080 8200 5082
rect 8412 5080 8458 5082
rect 1820 5067 2040 5080
rect 5832 5070 6060 5080
rect 6120 5070 6136 5080
rect 1818 5061 2040 5067
rect 1818 5060 1830 5061
rect 1800 5027 1830 5060
rect 1998 5027 2040 5061
rect 1800 4963 2040 5027
rect 2198 5061 2390 5067
rect 2198 5027 2210 5061
rect 2378 5027 2390 5061
rect 2198 5021 2390 5027
rect 2578 5061 3570 5067
rect 2578 5027 2590 5061
rect 3558 5027 3570 5061
rect 3758 5061 3950 5067
rect 3758 5040 3770 5061
rect 2578 5021 3570 5027
rect 3720 5027 3770 5040
rect 3938 5060 3950 5061
rect 3938 5027 3980 5060
rect 2142 4968 2188 4980
rect 1762 4960 2066 4963
rect 2142 4960 2148 4968
rect 1590 4840 1600 4960
rect 1720 4951 2148 4960
rect 1720 4840 1768 4951
rect 1762 4763 1768 4840
rect 1802 4840 2026 4951
rect 1802 4763 1808 4840
rect 1762 4751 1808 4763
rect 2020 4763 2026 4840
rect 2060 4840 2148 4951
rect 2060 4763 2066 4840
rect 2020 4751 2066 4763
rect 2142 4592 2148 4840
rect 2182 4960 2188 4968
rect 2400 4968 2446 4980
rect 2182 4840 2200 4960
rect 2182 4592 2188 4840
rect 2400 4800 2406 4968
rect 2440 4800 2446 4968
rect 2522 4968 2568 4980
rect 2142 4580 2188 4592
rect 2350 4580 2360 4800
rect 2440 4580 2450 4800
rect 2522 4760 2528 4968
rect 2520 4620 2528 4760
rect 2522 4592 2528 4620
rect 2562 4760 2568 4968
rect 3580 4968 3626 4980
rect 2562 4740 3380 4760
rect 2562 4620 3280 4740
rect 3380 4620 3390 4740
rect 2562 4592 2568 4620
rect 2522 4580 2568 4592
rect 3580 4592 3586 4968
rect 3620 4960 3626 4968
rect 3720 4963 3980 5027
rect 3702 4960 4006 4963
rect 3620 4951 4040 4960
rect 3620 4820 3708 4951
rect 3620 4592 3626 4820
rect 3702 4763 3708 4820
rect 3742 4820 3966 4951
rect 3742 4763 3748 4820
rect 3702 4751 3748 4763
rect 3960 4763 3966 4820
rect 4000 4840 4040 4951
rect 4140 4840 4150 4960
rect 5832 4894 5838 5070
rect 5872 4894 6060 5070
rect 6130 4894 6136 5070
rect 5832 4882 6060 4894
rect 5860 4880 6060 4882
rect 6120 4882 6136 4894
rect 6120 4880 6130 4882
rect 6330 4880 6340 5080
rect 6400 4880 6410 5080
rect 6570 4880 6580 5080
rect 6640 5070 6652 5080
rect 6646 4894 6652 5070
rect 6640 4882 6652 4894
rect 6640 4880 6650 4882
rect 6850 4880 6860 5080
rect 6920 4880 6930 5080
rect 7090 4880 7100 5080
rect 7160 5070 7170 5080
rect 7162 4894 7170 5070
rect 7160 4880 7170 4894
rect 7350 4880 7360 5080
rect 7420 4880 7430 5080
rect 7610 4880 7620 5080
rect 7680 4880 7690 5080
rect 7870 4880 7880 5080
rect 7940 4880 7950 5080
rect 8130 4880 8140 5080
rect 8200 4880 8210 5080
rect 8390 4880 8400 5080
rect 8460 4880 8470 5080
rect 8670 5070 8716 5082
rect 8928 5080 8974 5082
rect 9186 5080 9232 5082
rect 9444 5080 9490 5082
rect 9702 5080 9748 5082
rect 9960 5080 10006 5082
rect 10218 5080 10264 5082
rect 10476 5080 10522 5082
rect 10734 5080 10780 5082
rect 8650 4890 8660 5070
rect 8720 4890 8730 5070
rect 8670 4882 8716 4890
rect 8910 4880 8920 5080
rect 8980 4880 8990 5080
rect 9150 4880 9160 5080
rect 9220 5070 9232 5080
rect 9226 4894 9232 5070
rect 9220 4882 9232 4894
rect 9220 4880 9230 4882
rect 9410 4880 9420 5080
rect 9480 5070 9490 5080
rect 9484 4894 9490 5070
rect 9480 4880 9490 4894
rect 9670 4880 9680 5080
rect 9740 5070 9750 5080
rect 9742 4894 9750 5070
rect 9740 4880 9750 4894
rect 9930 4880 9940 5080
rect 10000 4880 10010 5080
rect 10190 4880 10200 5080
rect 10260 4880 10270 5080
rect 10450 4880 10460 5080
rect 10520 4880 10530 5080
rect 10710 5070 10780 5080
rect 10992 5070 11038 5082
rect 10710 4880 10720 5070
rect 10780 4880 10790 5070
rect 10992 5060 10998 5070
rect 11032 5060 11038 5070
rect 11250 5080 11554 5082
rect 11250 5070 11560 5080
rect 11250 5060 11256 5070
rect 11290 5060 11514 5070
rect 10970 4880 10980 5060
rect 11040 4880 11050 5060
rect 11230 4880 11240 5060
rect 11300 4894 11514 5060
rect 11548 4900 11560 5070
rect 11548 4894 11554 4900
rect 11300 4882 11554 4894
rect 11300 4880 11520 4882
rect 5860 4840 6100 4880
rect 6170 4840 6180 4860
rect 4000 4820 4020 4840
rect 4000 4763 4006 4820
rect 5860 4800 5900 4840
rect 6060 4800 6100 4840
rect 6160 4800 6180 4840
rect 6240 4840 6250 4860
rect 9550 4846 9630 4860
rect 6408 4840 6592 4846
rect 6668 4840 6852 4846
rect 7428 4840 7612 4846
rect 7688 4840 7872 4846
rect 8468 4840 8652 4846
rect 8728 4840 8912 4846
rect 9508 4840 9692 4846
rect 9748 4840 9932 4846
rect 10528 4840 10712 4846
rect 10788 4840 10972 4846
rect 11280 4840 11520 4880
rect 6240 4800 6420 4840
rect 6580 4800 6680 4840
rect 6840 4800 7440 4840
rect 7600 4800 7700 4840
rect 7860 4800 8480 4840
rect 8640 4800 8740 4840
rect 8900 4800 9520 4840
rect 9680 4800 9760 4840
rect 9920 4800 10540 4840
rect 10700 4800 10800 4840
rect 10960 4800 11220 4840
rect 11280 4800 11320 4840
rect 11480 4800 11520 4840
rect 5888 4794 6072 4800
rect 6408 4794 6592 4800
rect 6668 4794 6852 4800
rect 7428 4794 7612 4800
rect 7688 4794 7872 4800
rect 8468 4794 8652 4800
rect 8728 4794 8912 4800
rect 9508 4794 9692 4800
rect 9748 4794 9932 4800
rect 10528 4794 10712 4800
rect 10788 4794 10972 4800
rect 11308 4794 11492 4800
rect 3960 4751 4006 4763
rect 6560 4700 6580 4760
rect 6640 4700 7620 4760
rect 7680 4700 8660 4760
rect 8720 4700 9680 4760
rect 9740 4700 10720 4760
rect 10780 4700 10790 4760
rect 3580 4580 3626 4592
rect 4680 4640 5840 4660
rect 2200 4539 2620 4540
rect 1818 4533 2010 4539
rect 1818 4499 1830 4533
rect 1998 4499 2010 4533
rect 1818 4493 2010 4499
rect 2198 4533 2620 4539
rect 2720 4539 2730 4540
rect 2720 4533 3570 4539
rect 2198 4499 2210 4533
rect 2378 4500 2590 4533
rect 2378 4499 2390 4500
rect 2198 4493 2390 4499
rect 2578 4499 2590 4500
rect 3558 4499 3570 4533
rect 2578 4493 2620 4499
rect 2610 4480 2620 4493
rect 2720 4493 3570 4499
rect 3758 4533 3950 4539
rect 3758 4499 3770 4533
rect 3938 4499 3950 4533
rect 3758 4493 3950 4499
rect 2720 4480 2730 4493
rect 4680 4480 4700 4640
rect 4880 4600 5840 4640
rect 4880 4540 6180 4600
rect 6240 4540 6250 4600
rect 4880 4480 5840 4540
rect 6810 4500 6820 4560
rect 6880 4500 7220 4560
rect 7280 4500 7880 4560
rect 7940 4500 8900 4560
rect 8960 4500 9940 4560
rect 10000 4500 10960 4560
rect 11020 4500 12000 4560
rect 12060 4500 12070 4560
rect 4680 4460 5840 4480
rect 438 4381 630 4387
rect 438 4347 450 4381
rect 618 4380 630 4381
rect 818 4381 1010 4387
rect 618 4347 640 4380
rect 438 4341 640 4347
rect 818 4347 830 4381
rect 998 4347 1010 4381
rect 818 4341 1010 4347
rect 1076 4381 1268 4387
rect 1076 4347 1088 4381
rect 1256 4347 1268 4381
rect 1076 4341 1268 4347
rect 1458 4381 1650 4387
rect 1458 4347 1470 4381
rect 1638 4347 1650 4381
rect 1458 4341 1650 4347
rect 1716 4381 1908 4387
rect 1716 4347 1728 4381
rect 1896 4347 1908 4381
rect 1716 4341 1908 4347
rect 1974 4381 2166 4387
rect 1974 4347 1986 4381
rect 2154 4347 2166 4381
rect 1974 4341 2166 4347
rect 2232 4381 2424 4387
rect 2232 4347 2244 4381
rect 2412 4347 2424 4381
rect 2232 4341 2424 4347
rect 2618 4381 2810 4387
rect 2618 4347 2630 4381
rect 2798 4347 2810 4381
rect 2618 4341 2810 4347
rect 2876 4381 3068 4387
rect 2876 4347 2888 4381
rect 3056 4347 3068 4381
rect 2876 4341 3068 4347
rect 3134 4381 3326 4387
rect 3134 4347 3146 4381
rect 3314 4347 3326 4381
rect 3134 4341 3326 4347
rect 3392 4381 3584 4387
rect 3392 4347 3404 4381
rect 3572 4347 3584 4381
rect 3392 4341 3584 4347
rect 3778 4381 3970 4387
rect 3778 4347 3790 4381
rect 3958 4347 3970 4381
rect 7350 4380 7360 4440
rect 7420 4380 8400 4440
rect 8460 4380 9420 4440
rect 9480 4380 10440 4440
rect 10500 4380 10600 4440
rect 10660 4380 11480 4440
rect 11540 4380 11600 4440
rect 11660 4380 11670 4440
rect 14500 4403 14620 4420
rect 3778 4341 3970 4347
rect 440 4300 640 4341
rect 14500 4340 14566 4403
rect 5982 4320 6174 4326
rect 310 4220 320 4300
rect 400 4283 1060 4300
rect 400 4271 1066 4283
rect 422 4220 646 4271
rect 382 4083 388 4220
rect 422 4083 428 4220
rect 382 4071 428 4083
rect 640 4083 646 4220
rect 680 4220 1026 4271
rect 680 4083 686 4220
rect 640 4071 686 4083
rect 762 4117 808 4129
rect 762 4020 768 4117
rect 760 3929 768 4020
rect 802 4020 808 4117
rect 1020 4083 1026 4220
rect 1060 4083 1066 4271
rect 1660 4271 2360 4300
rect 1020 4071 1066 4083
rect 1278 4117 1324 4129
rect 1278 4020 1284 4117
rect 802 3929 1284 4020
rect 1318 3929 1324 4117
rect 1402 4117 1448 4129
rect 1402 4000 1408 4117
rect 760 3917 1324 3929
rect 1400 3929 1408 4000
rect 1442 4000 1448 4117
rect 1660 4083 1666 4271
rect 1700 4200 2182 4271
rect 1700 4083 1706 4200
rect 1660 4071 1706 4083
rect 1918 4117 1964 4129
rect 1918 4000 1924 4117
rect 1442 3929 1924 4000
rect 1958 4000 1964 4117
rect 2176 4083 2182 4200
rect 2216 4200 2360 4271
rect 2440 4200 2500 4300
rect 5960 4286 5994 4320
rect 6162 4286 6174 4320
rect 2820 4280 2866 4283
rect 3336 4280 3382 4283
rect 2820 4271 2920 4280
rect 2216 4083 2222 4200
rect 2176 4071 2222 4083
rect 2434 4117 2480 4129
rect 2434 4000 2440 4117
rect 1958 3929 2440 4000
rect 2474 4000 2480 4117
rect 2562 4117 2608 4129
rect 2562 4000 2568 4117
rect 2474 3929 2568 4000
rect 2602 4000 2608 4117
rect 2820 4083 2826 4271
rect 2860 4180 2920 4271
rect 3020 4271 3382 4280
rect 3020 4180 3342 4271
rect 2860 4083 2866 4180
rect 2820 4071 2866 4083
rect 3078 4117 3124 4129
rect 3078 4000 3084 4117
rect 2602 3929 3084 4000
rect 3118 4000 3124 4117
rect 3336 4083 3342 4180
rect 3376 4083 3382 4271
rect 5960 4280 6174 4286
rect 6240 4320 6432 4326
rect 6240 4286 6252 4320
rect 6420 4286 6432 4320
rect 6240 4280 6432 4286
rect 6498 4320 6690 4326
rect 6498 4286 6510 4320
rect 6678 4286 6690 4320
rect 6498 4280 6690 4286
rect 6902 4320 7094 4326
rect 6902 4286 6914 4320
rect 7082 4286 7094 4320
rect 6902 4280 7094 4286
rect 7160 4320 7352 4326
rect 7160 4286 7172 4320
rect 7340 4286 7352 4320
rect 7160 4280 7352 4286
rect 7418 4320 7610 4326
rect 7418 4286 7430 4320
rect 7598 4286 7610 4320
rect 7418 4280 7610 4286
rect 7676 4320 7868 4326
rect 7676 4286 7688 4320
rect 7856 4286 7868 4320
rect 7676 4280 7868 4286
rect 7934 4320 8126 4326
rect 7934 4286 7946 4320
rect 8114 4286 8126 4320
rect 7934 4280 8126 4286
rect 8192 4320 8384 4326
rect 8192 4286 8204 4320
rect 8372 4286 8384 4320
rect 8192 4280 8384 4286
rect 8450 4320 8642 4326
rect 8450 4286 8462 4320
rect 8630 4286 8642 4320
rect 8450 4280 8642 4286
rect 8708 4320 8900 4326
rect 8708 4286 8720 4320
rect 8888 4286 8900 4320
rect 8708 4280 8900 4286
rect 8966 4320 9158 4326
rect 8966 4286 8978 4320
rect 9146 4286 9158 4320
rect 8966 4280 9158 4286
rect 9224 4320 9416 4326
rect 9224 4286 9236 4320
rect 9404 4286 9416 4320
rect 9224 4280 9416 4286
rect 9482 4320 9674 4326
rect 9482 4286 9494 4320
rect 9662 4286 9674 4320
rect 9482 4280 9674 4286
rect 9740 4320 9932 4326
rect 9740 4286 9752 4320
rect 9920 4286 9932 4320
rect 9740 4280 9932 4286
rect 9998 4320 10190 4326
rect 9998 4286 10010 4320
rect 10178 4286 10190 4320
rect 9998 4280 10190 4286
rect 10256 4320 10448 4326
rect 10256 4286 10268 4320
rect 10436 4286 10448 4320
rect 10256 4280 10448 4286
rect 10514 4320 10706 4326
rect 10514 4286 10526 4320
rect 10694 4286 10706 4320
rect 10514 4280 10706 4286
rect 10772 4320 10964 4326
rect 10772 4286 10784 4320
rect 10952 4286 10964 4320
rect 10772 4280 10964 4286
rect 11030 4320 11222 4326
rect 11030 4286 11042 4320
rect 11210 4286 11222 4320
rect 11030 4280 11222 4286
rect 11288 4320 11480 4326
rect 11288 4286 11300 4320
rect 11468 4286 11480 4320
rect 11288 4280 11480 4286
rect 11546 4320 11738 4326
rect 11546 4286 11558 4320
rect 11726 4286 11738 4320
rect 11546 4280 11738 4286
rect 11804 4320 11996 4326
rect 11804 4286 11816 4320
rect 11984 4286 11996 4320
rect 11804 4280 11996 4286
rect 12062 4320 12254 4326
rect 14300 4320 14566 4340
rect 12062 4286 12074 4320
rect 12242 4286 12320 4320
rect 12062 4280 12320 4286
rect 5960 4248 6140 4280
rect 5926 4240 6140 4248
rect 6184 4240 6230 4248
rect 5926 4236 6180 4240
rect 3336 4071 3382 4083
rect 3594 4117 3640 4129
rect 3594 4000 3600 4117
rect 3118 3929 3600 4000
rect 3634 4000 3640 4117
rect 3722 4117 3768 4129
rect 3722 4000 3728 4117
rect 3634 3929 3728 4000
rect 3762 4000 3768 4117
rect 3980 4117 4026 4129
rect 3980 4000 3986 4117
rect 3762 3929 3986 4000
rect 4020 4000 4026 4117
rect 5926 4060 5932 4236
rect 5966 4080 6180 4236
rect 5966 4060 6140 4080
rect 6170 4060 6180 4080
rect 6240 4100 6250 4240
rect 6442 4236 6488 4248
rect 6442 4200 6448 4236
rect 6482 4200 6488 4236
rect 6700 4240 6746 4248
rect 6700 4236 6800 4240
rect 6700 4200 6706 4236
rect 6740 4200 6800 4236
rect 6846 4236 6892 4248
rect 6846 4220 6852 4236
rect 6886 4220 6892 4236
rect 7104 4236 7150 4248
rect 7104 4220 7110 4236
rect 7144 4220 7150 4236
rect 7362 4236 7408 4248
rect 7362 4220 7368 4236
rect 7402 4220 7408 4236
rect 7620 4236 7666 4248
rect 7620 4220 7626 4236
rect 7660 4220 7666 4236
rect 7878 4236 7924 4248
rect 7878 4220 7884 4236
rect 7918 4220 7924 4236
rect 8136 4236 8182 4248
rect 8136 4220 8142 4236
rect 8176 4220 8182 4236
rect 8394 4236 8440 4248
rect 8394 4220 8400 4236
rect 8434 4220 8440 4236
rect 8652 4236 8698 4248
rect 8652 4220 8658 4236
rect 8692 4220 8698 4236
rect 8910 4236 8956 4248
rect 8910 4220 8916 4236
rect 8950 4220 8956 4236
rect 9168 4236 9214 4248
rect 9168 4220 9174 4236
rect 9208 4220 9214 4236
rect 9426 4236 9472 4248
rect 9426 4220 9432 4236
rect 9466 4220 9472 4236
rect 9684 4236 9730 4248
rect 9684 4220 9690 4236
rect 9724 4220 9730 4236
rect 9942 4236 9988 4248
rect 9942 4220 9948 4236
rect 9982 4220 9988 4236
rect 10200 4236 10246 4248
rect 10200 4220 10206 4236
rect 10240 4220 10246 4236
rect 10458 4236 10504 4248
rect 10458 4220 10464 4236
rect 10498 4220 10504 4236
rect 10716 4236 10762 4248
rect 10716 4220 10722 4236
rect 10756 4220 10762 4236
rect 10974 4236 11020 4248
rect 10974 4220 10980 4236
rect 11014 4220 11020 4236
rect 11232 4236 11278 4248
rect 11232 4220 11238 4236
rect 11272 4220 11278 4236
rect 11490 4236 11536 4248
rect 11490 4220 11496 4236
rect 11530 4220 11536 4236
rect 11748 4236 11794 4248
rect 11748 4220 11754 4236
rect 11788 4220 11794 4236
rect 12006 4236 12052 4248
rect 12006 4220 12012 4236
rect 12046 4220 12052 4236
rect 12100 4236 12320 4280
rect 12100 4220 12270 4236
rect 6240 4060 6320 4100
rect 6430 4060 6440 4200
rect 6500 4060 6510 4200
rect 6690 4060 6700 4200
rect 6760 4080 6800 4200
rect 6760 4060 6770 4080
rect 6830 4060 6840 4220
rect 6900 4120 6910 4220
rect 6900 4060 6960 4120
rect 7090 4060 7100 4220
rect 7160 4060 7170 4220
rect 7350 4060 7360 4220
rect 7420 4060 7430 4220
rect 7610 4060 7620 4220
rect 7680 4060 7690 4220
rect 7870 4060 7880 4220
rect 7940 4060 7950 4220
rect 8130 4060 8140 4220
rect 8200 4060 8210 4220
rect 8390 4060 8400 4220
rect 8460 4060 8470 4220
rect 8630 4060 8640 4220
rect 8700 4060 8710 4220
rect 8890 4060 8900 4220
rect 8960 4060 8970 4220
rect 9150 4060 9160 4220
rect 9220 4060 9230 4220
rect 9410 4060 9420 4220
rect 9480 4060 9490 4220
rect 9670 4060 9680 4220
rect 9740 4060 9750 4220
rect 9930 4060 9940 4220
rect 10000 4060 10010 4220
rect 10190 4060 10200 4220
rect 10260 4060 10270 4220
rect 10430 4060 10440 4220
rect 10500 4060 10530 4220
rect 10690 4060 10700 4220
rect 10760 4060 10790 4220
rect 10950 4060 10960 4220
rect 11020 4060 11030 4220
rect 11210 4060 11220 4220
rect 11280 4060 11290 4220
rect 11470 4060 11480 4220
rect 11540 4060 11550 4220
rect 11730 4060 11740 4220
rect 11800 4060 11810 4220
rect 11990 4060 12000 4220
rect 12060 4080 12270 4220
rect 12060 4060 12070 4080
rect 12100 4060 12270 4080
rect 12304 4060 12320 4236
rect 14300 4160 14320 4320
rect 14460 4160 14566 4320
rect 14300 4140 14566 4160
rect 5926 4048 6140 4060
rect 6184 4048 6320 4060
rect 6442 4048 6488 4060
rect 6700 4048 6746 4060
rect 6846 4048 6960 4060
rect 7104 4048 7150 4060
rect 7362 4048 7408 4060
rect 7620 4048 7666 4060
rect 7878 4048 7924 4060
rect 8136 4048 8182 4060
rect 8394 4048 8440 4060
rect 8652 4048 8698 4060
rect 8910 4048 8956 4060
rect 9168 4048 9214 4060
rect 9426 4048 9472 4060
rect 9684 4048 9730 4060
rect 9942 4048 9988 4060
rect 10200 4048 10246 4060
rect 10458 4048 10504 4060
rect 10716 4048 10762 4060
rect 10974 4048 11020 4060
rect 11232 4048 11278 4060
rect 11490 4048 11536 4060
rect 11748 4048 11794 4060
rect 12006 4048 12052 4060
rect 5960 4016 6140 4048
rect 6220 4020 6320 4048
rect 6860 4020 6960 4048
rect 6220 4016 6680 4020
rect 6860 4016 11960 4020
rect 12100 4016 12320 4060
rect 5960 4010 6174 4016
rect 4020 3929 4040 4000
rect 5960 3980 5994 4010
rect 5982 3976 5994 3980
rect 6162 3976 6174 4010
rect 6220 4010 6690 4016
rect 6220 4000 6252 4010
rect 5982 3970 6174 3976
rect 6240 3976 6252 4000
rect 6420 3980 6510 4010
rect 6420 3976 6432 3980
rect 6240 3970 6432 3976
rect 6498 3976 6510 3980
rect 6678 3976 6690 4010
rect 6860 4010 11996 4016
rect 6860 3980 6914 4010
rect 6498 3970 6690 3976
rect 6902 3976 6914 3980
rect 7082 3980 7172 4010
rect 7082 3976 7094 3980
rect 6902 3970 7094 3976
rect 7160 3976 7172 3980
rect 7340 3980 7430 4010
rect 7340 3976 7352 3980
rect 7160 3970 7352 3976
rect 7418 3976 7430 3980
rect 7598 3980 7688 4010
rect 7598 3976 7610 3980
rect 7418 3970 7610 3976
rect 7676 3976 7688 3980
rect 7856 3980 7946 4010
rect 7856 3976 7868 3980
rect 7676 3970 7868 3976
rect 7934 3976 7946 3980
rect 8114 3980 8204 4010
rect 8114 3976 8126 3980
rect 7934 3970 8126 3976
rect 8192 3976 8204 3980
rect 8372 3980 8462 4010
rect 8372 3976 8384 3980
rect 8192 3970 8384 3976
rect 8450 3976 8462 3980
rect 8630 3980 8720 4010
rect 8630 3976 8642 3980
rect 8450 3970 8642 3976
rect 8708 3976 8720 3980
rect 8888 3980 8978 4010
rect 8888 3976 8900 3980
rect 8708 3970 8900 3976
rect 8966 3976 8978 3980
rect 9146 3980 9236 4010
rect 9146 3976 9158 3980
rect 8966 3970 9158 3976
rect 9224 3976 9236 3980
rect 9404 3980 9494 4010
rect 9404 3976 9416 3980
rect 9224 3970 9416 3976
rect 9482 3976 9494 3980
rect 9662 3980 9752 4010
rect 9662 3976 9674 3980
rect 9482 3970 9674 3976
rect 9740 3976 9752 3980
rect 9920 3980 10010 4010
rect 9920 3976 9932 3980
rect 9740 3970 9932 3976
rect 9998 3976 10010 3980
rect 10178 3980 10268 4010
rect 10178 3976 10190 3980
rect 9998 3970 10190 3976
rect 10256 3976 10268 3980
rect 10436 3980 10526 4010
rect 10436 3976 10448 3980
rect 10256 3970 10448 3976
rect 10514 3976 10526 3980
rect 10694 3980 10784 4010
rect 10694 3976 10706 3980
rect 10514 3970 10706 3976
rect 10772 3976 10784 3980
rect 10952 3980 11042 4010
rect 10952 3976 10964 3980
rect 10772 3970 10964 3976
rect 11030 3976 11042 3980
rect 11210 3980 11300 4010
rect 11210 3976 11222 3980
rect 11030 3970 11222 3976
rect 11288 3976 11300 3980
rect 11468 3980 11558 4010
rect 11468 3976 11480 3980
rect 11288 3970 11480 3976
rect 11546 3976 11558 3980
rect 11726 3980 11816 4010
rect 11726 3976 11738 3980
rect 11546 3970 11738 3976
rect 11804 3976 11816 3980
rect 11984 3976 11996 4010
rect 11804 3970 11996 3976
rect 12062 4010 12320 4016
rect 12062 3976 12074 4010
rect 12242 3980 12320 4010
rect 14500 4006 14566 4140
rect 14604 4006 14620 4403
rect 14726 4403 14776 4415
rect 14726 4400 14732 4403
rect 14500 4000 14620 4006
rect 14720 4006 14732 4400
rect 14770 4400 14776 4403
rect 14892 4403 14942 4415
rect 14892 4400 14898 4403
rect 14770 4006 14898 4400
rect 14936 4006 14942 4403
rect 14720 4000 14942 4006
rect 14560 3994 14610 4000
rect 14726 3994 14776 4000
rect 14892 3994 14942 4000
rect 15058 4403 15108 4415
rect 15058 4006 15064 4403
rect 15102 4400 15108 4403
rect 15224 4403 15274 4415
rect 15224 4400 15230 4403
rect 15102 4006 15230 4400
rect 15268 4400 15274 4403
rect 15390 4403 15440 4415
rect 15390 4400 15396 4403
rect 15268 4006 15280 4400
rect 15058 4000 15280 4006
rect 15380 4006 15396 4400
rect 15434 4400 15440 4403
rect 15556 4403 15606 4415
rect 15556 4400 15562 4403
rect 15434 4006 15562 4400
rect 15600 4006 15606 4403
rect 15380 4000 15606 4006
rect 15058 3994 15108 4000
rect 15224 3994 15274 4000
rect 15390 3994 15440 4000
rect 15556 3994 15606 4000
rect 15722 4403 15772 4415
rect 15722 4006 15728 4403
rect 15766 4400 15772 4403
rect 16034 4403 16084 4415
rect 16034 4400 16040 4403
rect 15766 4380 16040 4400
rect 15766 4020 15860 4380
rect 15940 4020 16040 4380
rect 15766 4006 16040 4020
rect 16078 4006 16084 4403
rect 15722 4000 16084 4006
rect 15722 3994 15772 4000
rect 16034 3994 16084 4000
rect 16200 4403 16250 4415
rect 16200 4006 16206 4403
rect 16244 4400 16250 4403
rect 16366 4403 16416 4415
rect 16366 4400 16372 4403
rect 16244 4006 16372 4400
rect 16410 4400 16416 4403
rect 16532 4403 16582 4415
rect 16410 4006 16440 4400
rect 16200 4000 16440 4006
rect 16532 4006 16538 4403
rect 16576 4400 16582 4403
rect 16698 4403 16748 4415
rect 16698 4400 16704 4403
rect 16576 4006 16704 4400
rect 16742 4400 16748 4403
rect 16864 4403 16914 4415
rect 16864 4400 16870 4403
rect 16742 4006 16760 4400
rect 16532 4000 16760 4006
rect 16860 4006 16870 4400
rect 16908 4400 16914 4403
rect 17030 4403 17080 4415
rect 17030 4400 17036 4403
rect 16908 4006 17036 4400
rect 17074 4006 17080 4403
rect 17196 4403 17246 4415
rect 17196 4040 17202 4403
rect 16860 4000 17080 4006
rect 16200 3994 16250 4000
rect 16366 3994 16416 4000
rect 16532 3994 16582 4000
rect 16698 3994 16748 4000
rect 16864 3994 16914 4000
rect 17030 3994 17080 4000
rect 17180 4006 17202 4040
rect 17240 4040 17246 4403
rect 17240 4006 17260 4040
rect 12242 3976 12254 3980
rect 12062 3970 12254 3976
rect 17180 3960 17260 4006
rect 760 3860 1320 3917
rect 1400 3900 4040 3929
rect 16760 3940 17260 3960
rect 6028 3920 6392 3926
rect 6028 3900 6040 3920
rect 438 3853 630 3859
rect 438 3819 450 3853
rect 618 3819 630 3853
rect 760 3853 840 3860
rect 940 3859 2420 3860
rect 940 3853 2424 3859
rect 760 3840 830 3853
rect 438 3813 630 3819
rect 818 3819 830 3840
rect 998 3819 1088 3853
rect 1256 3819 1470 3853
rect 1638 3819 1728 3853
rect 1896 3819 1986 3853
rect 2154 3819 2244 3853
rect 2412 3819 2424 3853
rect 818 3813 840 3819
rect 820 3800 840 3813
rect 940 3813 2424 3819
rect 940 3800 2420 3813
rect 2610 3800 2620 3860
rect 2720 3859 3580 3860
rect 3780 3859 3960 3900
rect 2720 3853 3584 3859
rect 2798 3820 2888 3853
rect 2798 3819 2810 3820
rect 2720 3813 2810 3819
rect 2876 3819 2888 3820
rect 3056 3820 3146 3853
rect 3056 3819 3068 3820
rect 2876 3813 3068 3819
rect 3134 3819 3146 3820
rect 3314 3820 3404 3853
rect 3314 3819 3326 3820
rect 3134 3813 3326 3819
rect 3392 3819 3404 3820
rect 3572 3819 3584 3853
rect 3392 3813 3584 3819
rect 3778 3853 3970 3859
rect 3778 3819 3790 3853
rect 3958 3819 3970 3853
rect 3778 3813 3970 3819
rect 2720 3800 2730 3813
rect 5640 3700 5660 3900
rect 5840 3860 6040 3900
rect 6380 3900 6392 3920
rect 6380 3860 6440 3900
rect 5840 3840 6440 3860
rect 6500 3840 7100 3900
rect 7160 3840 7620 3900
rect 7680 3840 8140 3900
rect 8200 3840 8640 3900
rect 8700 3840 9160 3900
rect 9220 3840 9680 3900
rect 9740 3840 10200 3900
rect 10260 3840 10700 3900
rect 10760 3840 11220 3900
rect 11280 3840 11740 3900
rect 11800 3840 12070 3900
rect 16760 3880 16780 3940
rect 16860 3880 17260 3940
rect 5840 3700 6380 3840
rect 17170 3800 17180 3820
rect 15850 3720 15860 3800
rect 15940 3720 17180 3800
rect 17260 3720 17270 3820
rect 15860 3700 17260 3720
rect 4040 3540 4370 3560
rect 2610 3420 2620 3540
rect 2720 3420 4370 3540
rect 17170 3460 17180 3520
rect 17240 3500 17250 3520
rect 17240 3494 17260 3500
rect 17242 3460 17260 3494
rect 17196 3454 17254 3460
rect 2620 3400 4370 3420
rect 4040 3360 4370 3400
rect 12870 3240 12880 3440
rect 13080 3370 14500 3440
rect 13080 3260 16900 3370
rect 16970 3260 16980 3370
rect 13080 3240 14500 3260
rect 380 3141 640 3160
rect 380 3107 430 3141
rect 598 3107 640 3141
rect 380 3043 640 3107
rect 798 3141 990 3147
rect 798 3107 810 3141
rect 978 3107 990 3141
rect 798 3101 990 3107
rect 1056 3141 1248 3147
rect 1056 3107 1068 3141
rect 1236 3107 1248 3141
rect 1056 3101 1248 3107
rect 1314 3141 1506 3147
rect 1314 3107 1326 3141
rect 1494 3107 1506 3141
rect 1314 3101 1506 3107
rect 1572 3141 1764 3147
rect 1572 3107 1584 3141
rect 1752 3107 1764 3141
rect 1572 3101 1764 3107
rect 1830 3141 2022 3147
rect 1830 3107 1842 3141
rect 2010 3107 2022 3141
rect 1830 3101 2022 3107
rect 2088 3141 2280 3147
rect 2088 3107 2100 3141
rect 2268 3107 2280 3141
rect 2088 3101 2280 3107
rect 2346 3141 2538 3147
rect 2346 3107 2358 3141
rect 2526 3107 2538 3141
rect 2346 3101 2538 3107
rect 2604 3141 2796 3147
rect 2604 3107 2616 3141
rect 2784 3107 2796 3141
rect 2604 3101 2796 3107
rect 2960 3141 3180 3160
rect 2960 3107 2990 3141
rect 3158 3107 3180 3141
rect 2960 3043 3180 3107
rect 362 3040 666 3043
rect 1000 3040 1046 3043
rect 1516 3040 1562 3043
rect 2032 3040 2078 3043
rect 2548 3040 2594 3043
rect 2922 3040 3226 3043
rect 3274 3040 3366 3052
rect 4040 3040 4380 3100
rect 360 3031 3280 3040
rect 360 2940 368 3031
rect 362 2843 368 2940
rect 402 2940 626 3031
rect 402 2843 408 2940
rect 362 2831 408 2843
rect 620 2843 626 2940
rect 660 2940 1006 3031
rect 660 2843 666 2940
rect 620 2831 666 2843
rect 742 2877 788 2889
rect 742 2800 748 2877
rect 740 2689 748 2800
rect 782 2800 788 2877
rect 1000 2843 1006 2940
rect 1040 2940 1522 3031
rect 1040 2843 1046 2940
rect 1000 2831 1046 2843
rect 1258 2877 1304 2889
rect 1258 2800 1264 2877
rect 782 2689 1264 2800
rect 1298 2800 1304 2877
rect 1516 2843 1522 2940
rect 1556 2940 2038 3031
rect 1556 2843 1562 2940
rect 1516 2831 1562 2843
rect 1774 2877 1820 2889
rect 1774 2800 1780 2877
rect 1298 2689 1780 2800
rect 1814 2800 1820 2877
rect 2032 2843 2038 2940
rect 2072 2940 2554 3031
rect 2072 2843 2078 2940
rect 2032 2831 2078 2843
rect 2290 2877 2336 2889
rect 2290 2800 2296 2877
rect 1814 2689 2296 2800
rect 2330 2800 2336 2877
rect 2548 2843 2554 2940
rect 2588 2940 2928 3031
rect 2588 2843 2594 2940
rect 2548 2831 2594 2843
rect 2806 2877 2852 2889
rect 2806 2800 2812 2877
rect 2330 2780 2812 2800
rect 2330 2689 2620 2780
rect 418 2613 610 2619
rect 418 2579 430 2613
rect 598 2579 610 2613
rect 418 2573 610 2579
rect 740 2613 2620 2689
rect 2700 2689 2812 2780
rect 2846 2689 2852 2877
rect 2922 2843 2928 2940
rect 2962 2940 3186 3031
rect 2962 2843 2968 2940
rect 2922 2831 2968 2843
rect 3180 2843 3186 2940
rect 3220 2940 3280 3031
rect 3400 2940 4380 3040
rect 3220 2843 3226 2940
rect 3274 2928 3366 2940
rect 4040 2900 4380 2940
rect 4560 2900 4580 3100
rect 14300 3080 14500 3120
rect 14300 2940 14340 3080
rect 14460 3060 14500 3080
rect 14460 3029 16714 3060
rect 14460 2995 14627 3029
rect 14661 2995 14719 3029
rect 14753 2995 14811 3029
rect 14845 2995 14903 3029
rect 14937 2995 14995 3029
rect 15029 2995 15087 3029
rect 15121 2995 15179 3029
rect 15213 2995 15271 3029
rect 15305 2995 15363 3029
rect 15397 2995 15455 3029
rect 15489 2995 15547 3029
rect 15581 2995 15639 3029
rect 15673 2995 15731 3029
rect 15765 2995 15823 3029
rect 15857 2995 15915 3029
rect 15949 2995 16007 3029
rect 16041 2995 16099 3029
rect 16133 2995 16191 3029
rect 16225 2995 16283 3029
rect 16317 2995 16375 3029
rect 16409 2995 16467 3029
rect 16501 2995 16559 3029
rect 16593 2995 16651 3029
rect 16685 2995 16714 3029
rect 14460 2964 16714 2995
rect 14460 2960 14640 2964
rect 14300 2920 14430 2940
rect 14420 2910 14430 2920
rect 14500 2910 14520 2960
rect 14420 2880 14520 2910
rect 3180 2831 3226 2843
rect 14789 2859 14847 2865
rect 14789 2825 14801 2859
rect 14835 2856 14847 2859
rect 15167 2859 15225 2865
rect 15167 2856 15179 2859
rect 14835 2828 15179 2856
rect 14835 2825 14847 2828
rect 14789 2819 14847 2825
rect 15167 2825 15179 2828
rect 15213 2856 15225 2859
rect 15791 2859 15849 2865
rect 15791 2856 15803 2859
rect 15213 2828 15803 2856
rect 15213 2825 15225 2828
rect 15167 2819 15225 2825
rect 15791 2825 15803 2828
rect 15837 2825 15849 2859
rect 17070 2840 17080 3420
rect 17140 3413 17180 3420
rect 17140 3401 17204 3413
rect 17140 2840 17164 3401
rect 15791 2819 15849 2825
rect 17158 2825 17164 2840
rect 17198 2825 17204 3401
rect 17158 2813 17204 2825
rect 17246 3401 17292 3413
rect 17246 2825 17252 3401
rect 17286 3400 17292 3401
rect 17354 3400 17406 3412
rect 17286 2840 17360 3400
rect 17400 3380 17440 3400
rect 17440 3300 17450 3380
rect 17400 3260 17440 3300
rect 17440 3180 17450 3260
rect 17400 3120 17440 3180
rect 17440 3040 17450 3120
rect 17400 2980 17440 3040
rect 17440 2900 17450 2980
rect 17400 2840 17440 2900
rect 17286 2825 17292 2840
rect 17354 2828 17406 2840
rect 17246 2813 17292 2825
rect 13080 2760 14500 2780
rect 17196 2766 17254 2772
rect 17196 2760 17208 2766
rect 17242 2760 17254 2766
rect 2700 2677 2852 2689
rect 2700 2613 2840 2677
rect 740 2579 810 2613
rect 978 2579 1068 2613
rect 1236 2579 1326 2613
rect 1494 2579 1584 2613
rect 1752 2579 1842 2613
rect 2010 2579 2100 2613
rect 2268 2579 2358 2613
rect 2526 2579 2616 2613
rect 2784 2579 2840 2613
rect 740 2560 2840 2579
rect 2978 2613 3170 2619
rect 2978 2579 2990 2613
rect 3158 2579 3170 2613
rect 13070 2580 13080 2760
rect 13260 2740 14500 2760
rect 14614 2740 14666 2752
rect 13260 2680 14620 2740
rect 14660 2680 14666 2740
rect 14708 2723 14766 2729
rect 14708 2689 14720 2723
rect 14754 2720 14766 2723
rect 15075 2723 15133 2729
rect 15075 2720 15087 2723
rect 14754 2692 15087 2720
rect 14754 2689 14766 2692
rect 14708 2683 14766 2689
rect 15075 2689 15087 2692
rect 15121 2720 15133 2723
rect 15791 2723 15849 2729
rect 15791 2720 15803 2723
rect 15121 2692 15803 2720
rect 15121 2689 15133 2692
rect 15075 2683 15133 2689
rect 15791 2689 15803 2692
rect 15837 2689 15849 2723
rect 15791 2683 15849 2689
rect 16007 2718 16065 2724
rect 16007 2684 16019 2718
rect 16053 2684 16065 2718
rect 13260 2580 14500 2680
rect 14614 2668 14666 2680
rect 16007 2661 16065 2684
rect 16638 2720 16702 2726
rect 16890 2720 16900 2740
rect 16638 2680 16650 2720
rect 16690 2680 16900 2720
rect 16638 2674 16702 2680
rect 15347 2660 15477 2661
rect 14880 2590 14890 2660
rect 14970 2590 14980 2660
rect 15330 2600 15340 2660
rect 15400 2655 15477 2660
rect 15400 2621 15431 2655
rect 15465 2652 15477 2655
rect 16007 2655 16125 2661
rect 16890 2660 16900 2680
rect 16980 2660 16990 2740
rect 17180 2720 17200 2760
rect 17190 2700 17200 2720
rect 17260 2700 17270 2760
rect 16007 2652 16079 2655
rect 15465 2624 16079 2652
rect 15465 2621 15477 2624
rect 15400 2615 15477 2621
rect 16067 2621 16079 2624
rect 16113 2621 16125 2655
rect 16067 2615 16125 2621
rect 16328 2620 16412 2626
rect 15400 2600 15410 2615
rect 2978 2573 3170 2579
rect 16328 2560 16340 2620
rect 16400 2560 16780 2620
rect 16860 2560 16870 2620
rect 16328 2554 16412 2560
rect 14598 2500 16714 2516
rect 2030 2420 2040 2480
rect 2100 2420 2920 2480
rect 3020 2420 3030 2480
rect 14598 2420 14620 2500
rect 14700 2485 16714 2500
rect 14700 2451 14719 2485
rect 14753 2451 14811 2485
rect 14845 2451 14903 2485
rect 14937 2451 14995 2485
rect 15029 2451 15087 2485
rect 15121 2451 15179 2485
rect 15213 2451 15271 2485
rect 15305 2451 15363 2485
rect 15397 2451 15455 2485
rect 15489 2451 15547 2485
rect 15581 2451 15639 2485
rect 15673 2451 15731 2485
rect 15765 2451 15823 2485
rect 15857 2451 15915 2485
rect 15949 2451 16007 2485
rect 16041 2451 16099 2485
rect 16133 2451 16191 2485
rect 16225 2451 16283 2485
rect 16317 2451 16375 2485
rect 16409 2451 16467 2485
rect 16501 2451 16559 2485
rect 16593 2451 16651 2485
rect 16685 2451 16714 2485
rect 14700 2420 16714 2451
rect 17190 2420 17200 2440
rect 17180 2380 17200 2420
rect 17260 2380 17270 2440
rect 530 2240 540 2320
rect 600 2300 1180 2320
rect 600 2240 840 2300
rect 940 2240 1180 2300
rect 1240 2240 1250 2320
rect 1290 2280 1300 2360
rect 1360 2280 1940 2360
rect 2000 2280 2620 2360
rect 2720 2280 2730 2360
rect 14890 2320 14900 2380
rect 14960 2370 17130 2380
rect 14960 2320 17060 2370
rect 17050 2310 17060 2320
rect 17120 2320 17130 2370
rect 17196 2372 17208 2380
rect 17242 2372 17254 2380
rect 17196 2366 17254 2372
rect 17158 2322 17204 2334
rect 17158 2320 17164 2322
rect 17120 2310 17164 2320
rect 14300 2200 14500 2220
rect 2690 2080 2700 2160
rect 2760 2080 2920 2160
rect 3000 2080 3010 2160
rect 14300 2020 14340 2200
rect 14460 2160 14500 2200
rect 14460 2100 15340 2160
rect 15400 2100 15410 2160
rect 17070 2146 17164 2310
rect 17198 2146 17204 2322
rect 17070 2140 17204 2146
rect 17158 2134 17204 2140
rect 17246 2322 17292 2334
rect 17246 2146 17252 2322
rect 17286 2320 17292 2322
rect 17286 2300 17460 2320
rect 17286 2280 17360 2300
rect 17400 2280 17460 2300
rect 17286 2146 17320 2280
rect 17246 2140 17320 2146
rect 17420 2140 17460 2280
rect 17246 2134 17292 2140
rect 17340 2120 17460 2140
rect 17196 2100 17254 2102
rect 14460 2020 14500 2100
rect 17180 2096 17260 2100
rect 17180 2062 17208 2096
rect 17242 2062 17260 2096
rect 17180 2060 17260 2062
rect 17196 2056 17254 2060
rect 160 1944 480 1970
rect 2670 1960 2680 1980
rect 160 1910 234 1944
rect 402 1910 480 1944
rect 600 1944 2680 1960
rect 600 1920 614 1944
rect 160 1860 480 1910
rect 602 1910 614 1920
rect 782 1920 994 1944
rect 782 1910 794 1920
rect 602 1904 794 1910
rect 982 1910 994 1920
rect 1162 1920 1374 1944
rect 1162 1910 1174 1920
rect 982 1904 1174 1910
rect 1362 1910 1374 1920
rect 1542 1920 1754 1944
rect 1542 1910 1554 1920
rect 1362 1904 1554 1910
rect 1742 1910 1754 1920
rect 1922 1920 2134 1944
rect 1922 1910 1934 1920
rect 1742 1904 1934 1910
rect 2122 1910 2134 1920
rect 2302 1920 2514 1944
rect 2760 1920 2770 1980
rect 2882 1944 3140 1950
rect 2882 1940 2894 1944
rect 2302 1910 2314 1920
rect 2122 1904 2314 1910
rect 2502 1910 2514 1920
rect 2682 1910 2694 1920
rect 2502 1904 2694 1910
rect 2860 1910 2894 1940
rect 3062 1910 3140 1944
rect 2860 1900 3140 1910
rect 546 1870 592 1872
rect 804 1870 850 1872
rect 926 1870 972 1872
rect 1184 1870 1230 1872
rect 160 1684 172 1860
rect 206 1684 430 1860
rect 464 1684 480 1860
rect 530 1690 540 1870
rect 600 1690 610 1870
rect 804 1860 820 1870
rect 960 1860 972 1870
rect 160 1634 480 1684
rect 546 1684 552 1690
rect 586 1684 592 1690
rect 546 1672 592 1684
rect 804 1684 810 1860
rect 966 1684 972 1860
rect 1170 1690 1180 1870
rect 1240 1690 1250 1870
rect 1306 1860 1352 1872
rect 1306 1850 1312 1860
rect 1346 1850 1352 1860
rect 1564 1870 1610 1872
rect 1686 1870 1732 1872
rect 1564 1860 1732 1870
rect 1944 1860 1990 1872
rect 2066 1870 2112 1872
rect 2324 1870 2370 1872
rect 2446 1870 2492 1872
rect 1290 1690 1300 1850
rect 1360 1690 1370 1850
rect 804 1672 820 1684
rect 810 1670 820 1672
rect 960 1672 972 1684
rect 1184 1684 1190 1690
rect 1224 1684 1230 1690
rect 1184 1672 1230 1684
rect 1306 1684 1312 1690
rect 1346 1684 1352 1690
rect 1306 1672 1352 1684
rect 1564 1684 1570 1860
rect 1604 1830 1692 1860
rect 1680 1690 1692 1830
rect 1604 1684 1692 1690
rect 1726 1684 1732 1860
rect 1564 1672 1732 1684
rect 1910 1680 1920 1860
rect 1984 1684 1990 1860
rect 1980 1680 1990 1684
rect 1944 1672 1990 1680
rect 960 1670 970 1672
rect 1580 1670 1720 1672
rect 2030 1670 2040 1870
rect 2120 1670 2130 1870
rect 2324 1860 2492 1870
rect 2324 1684 2330 1860
rect 2364 1850 2452 1860
rect 2364 1684 2370 1690
rect 2324 1672 2370 1684
rect 2446 1684 2452 1690
rect 2486 1684 2492 1860
rect 2704 1860 2750 1872
rect 2704 1850 2710 1860
rect 2446 1672 2492 1684
rect 2670 1670 2680 1850
rect 2744 1684 2750 1860
rect 2740 1670 2750 1684
rect 2820 1860 3140 1900
rect 2820 1684 2832 1860
rect 2866 1684 3090 1860
rect 3124 1684 3140 1860
rect 160 1600 234 1634
rect 402 1600 480 1634
rect 160 1526 480 1600
rect 602 1634 794 1640
rect 602 1600 614 1634
rect 782 1600 794 1634
rect 602 1594 794 1600
rect 982 1634 1174 1640
rect 982 1600 994 1634
rect 1162 1600 1174 1634
rect 982 1594 1174 1600
rect 1362 1634 1554 1640
rect 1362 1600 1374 1634
rect 1542 1600 1554 1634
rect 1362 1594 1554 1600
rect 1742 1634 1934 1640
rect 1742 1600 1754 1634
rect 1922 1600 1934 1634
rect 1742 1594 1934 1600
rect 2122 1634 2314 1640
rect 2122 1600 2134 1634
rect 2302 1600 2314 1634
rect 2122 1594 2314 1600
rect 2502 1634 2694 1640
rect 2502 1600 2514 1634
rect 2682 1600 2694 1634
rect 2502 1594 2694 1600
rect 2820 1634 3140 1684
rect 2820 1600 2894 1634
rect 3062 1600 3140 1634
rect 660 1532 760 1594
rect 1020 1532 1120 1594
rect 1400 1532 1500 1594
rect 1800 1532 1900 1594
rect 2180 1532 2280 1594
rect 2540 1532 2640 1594
rect 160 1492 234 1526
rect 402 1492 480 1526
rect 160 1442 480 1492
rect 602 1526 794 1532
rect 602 1492 614 1526
rect 782 1492 794 1526
rect 602 1486 794 1492
rect 982 1526 1174 1532
rect 982 1492 994 1526
rect 1162 1492 1174 1526
rect 982 1486 1174 1492
rect 1362 1526 1554 1532
rect 1362 1492 1374 1526
rect 1542 1492 1554 1526
rect 1362 1486 1554 1492
rect 1742 1526 1934 1532
rect 1742 1492 1754 1526
rect 1922 1492 1934 1526
rect 1742 1486 1934 1492
rect 2122 1526 2314 1532
rect 2122 1492 2134 1526
rect 2302 1492 2314 1526
rect 2122 1486 2314 1492
rect 2502 1526 2694 1532
rect 2502 1492 2514 1526
rect 2682 1492 2694 1526
rect 2502 1486 2694 1492
rect 2820 1526 3140 1600
rect 2820 1492 2894 1526
rect 3062 1492 3140 1526
rect 1020 1480 1120 1486
rect 1400 1480 1500 1486
rect 1800 1480 1900 1486
rect 2180 1480 2280 1486
rect 2540 1480 2640 1486
rect 546 1450 592 1454
rect 804 1450 850 1454
rect 926 1450 972 1454
rect 1184 1450 1230 1454
rect 160 1266 172 1442
rect 206 1266 430 1442
rect 464 1266 480 1442
rect 160 1216 480 1266
rect 530 1250 540 1450
rect 600 1250 610 1450
rect 804 1442 820 1450
rect 960 1442 972 1450
rect 804 1266 810 1442
rect 966 1266 972 1442
rect 1170 1270 1180 1450
rect 1240 1270 1250 1450
rect 1306 1442 1352 1454
rect 1306 1430 1312 1442
rect 1346 1430 1352 1442
rect 1564 1450 1610 1454
rect 1686 1450 1732 1454
rect 1564 1442 1732 1450
rect 1290 1270 1300 1430
rect 1360 1270 1370 1430
rect 804 1254 820 1266
rect 810 1250 820 1254
rect 960 1254 972 1266
rect 1184 1266 1190 1270
rect 1224 1266 1230 1270
rect 1184 1254 1230 1266
rect 1306 1266 1312 1270
rect 1346 1266 1352 1270
rect 1306 1254 1352 1266
rect 1564 1266 1570 1442
rect 1604 1410 1692 1442
rect 1604 1266 1692 1270
rect 1726 1266 1732 1442
rect 1944 1442 1990 1454
rect 2066 1450 2112 1454
rect 2324 1450 2370 1454
rect 2446 1450 2492 1454
rect 2704 1450 2750 1454
rect 1944 1440 1950 1442
rect 1564 1254 1732 1266
rect 1910 1260 1920 1440
rect 1984 1266 1990 1442
rect 1980 1260 1990 1266
rect 1944 1254 1990 1260
rect 960 1250 970 1254
rect 1580 1250 1720 1254
rect 2050 1250 2060 1450
rect 2140 1250 2150 1450
rect 2324 1442 2492 1450
rect 2324 1266 2330 1442
rect 2364 1430 2452 1442
rect 2364 1266 2370 1270
rect 2324 1254 2370 1266
rect 2446 1266 2452 1270
rect 2486 1266 2492 1442
rect 2690 1270 2700 1450
rect 2760 1270 2770 1450
rect 2820 1442 3140 1492
rect 2446 1254 2492 1266
rect 2704 1266 2710 1270
rect 2744 1266 2750 1270
rect 2704 1254 2750 1266
rect 2820 1266 2832 1442
rect 2866 1266 3090 1442
rect 3124 1266 3140 1442
rect 160 1182 234 1216
rect 402 1182 480 1216
rect 160 1108 480 1182
rect 602 1216 794 1222
rect 602 1182 614 1216
rect 782 1182 794 1216
rect 602 1176 794 1182
rect 982 1216 1174 1222
rect 982 1182 994 1216
rect 1162 1182 1174 1216
rect 982 1176 1174 1182
rect 1362 1216 1554 1222
rect 1362 1182 1374 1216
rect 1542 1182 1554 1216
rect 1362 1176 1554 1182
rect 1742 1216 1934 1222
rect 1742 1182 1754 1216
rect 1922 1182 1934 1216
rect 1742 1176 1934 1182
rect 2122 1216 2314 1222
rect 2122 1182 2134 1216
rect 2302 1182 2314 1216
rect 2122 1176 2314 1182
rect 2502 1216 2694 1222
rect 2502 1182 2514 1216
rect 2682 1182 2694 1216
rect 2502 1176 2694 1182
rect 2820 1216 3140 1266
rect 2820 1182 2894 1216
rect 3062 1182 3140 1216
rect 660 1114 760 1176
rect 1020 1114 1120 1176
rect 1400 1114 1500 1176
rect 1800 1114 1900 1176
rect 2180 1114 2280 1176
rect 2540 1114 2640 1176
rect 160 1074 234 1108
rect 402 1074 480 1108
rect 160 1024 480 1074
rect 602 1108 794 1114
rect 602 1074 614 1108
rect 782 1074 794 1108
rect 602 1068 794 1074
rect 982 1108 1174 1114
rect 982 1074 994 1108
rect 1162 1074 1174 1108
rect 982 1068 1174 1074
rect 1362 1108 1554 1114
rect 1362 1074 1374 1108
rect 1542 1074 1554 1108
rect 1362 1068 1554 1074
rect 1742 1108 1934 1114
rect 1742 1074 1754 1108
rect 1922 1074 1934 1108
rect 1742 1068 1934 1074
rect 2122 1108 2314 1114
rect 2122 1074 2134 1108
rect 2302 1074 2314 1108
rect 2122 1068 2314 1074
rect 2502 1108 2694 1114
rect 2502 1074 2514 1108
rect 2682 1074 2694 1108
rect 2502 1068 2694 1074
rect 2820 1108 3140 1182
rect 2820 1074 2894 1108
rect 3062 1074 3140 1108
rect 546 1030 592 1036
rect 804 1030 850 1036
rect 926 1030 972 1036
rect 1184 1030 1230 1036
rect 160 848 172 1024
rect 206 848 430 1024
rect 464 848 480 1024
rect 530 850 540 1030
rect 600 850 610 1030
rect 804 1024 820 1030
rect 960 1024 972 1030
rect 160 798 480 848
rect 546 848 552 850
rect 586 848 592 850
rect 546 836 592 848
rect 804 848 810 1024
rect 966 848 972 1024
rect 1170 850 1180 1030
rect 1240 850 1250 1030
rect 1306 1024 1352 1036
rect 1306 1010 1312 1024
rect 1346 1010 1352 1024
rect 1564 1030 1610 1036
rect 1686 1030 1732 1036
rect 1564 1024 1732 1030
rect 1290 850 1300 1010
rect 1360 850 1370 1010
rect 804 836 820 848
rect 810 830 820 836
rect 960 836 972 848
rect 1184 848 1190 850
rect 1224 848 1230 850
rect 1184 836 1230 848
rect 1306 848 1312 850
rect 1346 848 1352 850
rect 1306 836 1352 848
rect 1564 848 1570 1024
rect 1604 990 1692 1024
rect 1604 848 1692 850
rect 1726 848 1732 1024
rect 1944 1024 1990 1036
rect 2066 1030 2112 1036
rect 2324 1030 2370 1036
rect 2446 1030 2492 1036
rect 2704 1030 2750 1036
rect 1944 1020 1950 1024
rect 1564 836 1732 848
rect 1910 840 1920 1020
rect 1984 848 1990 1024
rect 2050 850 2060 1030
rect 2120 850 2130 1030
rect 2324 1024 2492 1030
rect 1980 840 1990 848
rect 1944 836 1990 840
rect 2066 848 2072 850
rect 2106 848 2112 850
rect 2066 836 2112 848
rect 2324 848 2330 1024
rect 2364 1010 2452 1024
rect 2364 848 2370 850
rect 2324 836 2370 848
rect 2446 848 2452 850
rect 2486 848 2492 1024
rect 2690 850 2700 1030
rect 2760 850 2770 1030
rect 2820 1024 3140 1074
rect 2446 836 2492 848
rect 2704 848 2710 850
rect 2744 848 2750 850
rect 2704 836 2750 848
rect 2820 848 2832 1024
rect 2866 848 3090 1024
rect 3124 848 3140 1024
rect 960 830 970 836
rect 1580 830 1720 836
rect 160 764 234 798
rect 402 764 480 798
rect 160 690 480 764
rect 602 798 794 804
rect 602 764 614 798
rect 782 764 794 798
rect 602 758 794 764
rect 982 798 1174 804
rect 982 764 994 798
rect 1162 764 1174 798
rect 982 758 1174 764
rect 1362 798 1554 804
rect 1362 764 1374 798
rect 1542 764 1554 798
rect 1362 758 1554 764
rect 1742 798 1934 804
rect 1742 764 1754 798
rect 1922 764 1934 798
rect 1742 758 1934 764
rect 2122 798 2314 804
rect 2122 764 2134 798
rect 2302 764 2314 798
rect 2122 758 2314 764
rect 2502 798 2694 804
rect 2502 764 2514 798
rect 2682 764 2694 798
rect 2502 758 2694 764
rect 2820 798 3140 848
rect 2820 764 2894 798
rect 3062 764 3140 798
rect 660 696 760 758
rect 1020 696 1120 758
rect 1400 696 1500 758
rect 1800 696 1900 758
rect 2180 696 2280 758
rect 2540 696 2640 758
rect 160 656 234 690
rect 402 656 480 690
rect 160 606 480 656
rect 602 690 794 696
rect 602 656 614 690
rect 782 656 794 690
rect 602 650 794 656
rect 982 690 1174 696
rect 982 656 994 690
rect 1162 656 1174 690
rect 982 650 1174 656
rect 1362 690 1554 696
rect 1362 656 1374 690
rect 1542 656 1554 690
rect 1362 650 1554 656
rect 1742 690 1934 696
rect 1742 656 1754 690
rect 1922 656 1934 690
rect 1742 650 1934 656
rect 2122 690 2314 696
rect 2122 656 2134 690
rect 2302 656 2314 690
rect 2122 650 2314 656
rect 2502 690 2694 696
rect 2502 656 2514 690
rect 2682 656 2694 690
rect 2502 650 2694 656
rect 2820 690 3140 764
rect 2820 656 2894 690
rect 3062 656 3140 690
rect 546 610 592 618
rect 804 610 850 618
rect 926 610 972 618
rect 1184 610 1230 618
rect 160 430 172 606
rect 206 430 430 606
rect 464 430 480 606
rect 530 430 540 610
rect 600 430 610 610
rect 804 606 820 610
rect 960 606 972 610
rect 804 430 810 606
rect 966 430 972 606
rect 1170 430 1180 610
rect 1240 430 1250 610
rect 1306 606 1352 618
rect 1306 590 1312 606
rect 1346 590 1352 606
rect 1564 610 1610 618
rect 1686 610 1732 618
rect 1564 606 1732 610
rect 1290 430 1300 590
rect 1360 430 1370 590
rect 1564 430 1570 606
rect 1604 570 1692 606
rect 1726 430 1732 606
rect 1944 606 1990 618
rect 2066 610 2112 618
rect 2324 610 2370 618
rect 2446 610 2492 618
rect 2704 610 2750 618
rect 1944 600 1950 606
rect 160 380 480 430
rect 546 418 592 430
rect 804 418 850 430
rect 926 418 972 430
rect 1184 418 1230 430
rect 1306 418 1352 430
rect 1564 418 1732 430
rect 1910 420 1920 600
rect 1984 430 1990 606
rect 2050 430 2060 610
rect 2120 430 2130 610
rect 2324 606 2492 610
rect 2324 430 2330 606
rect 2364 590 2452 606
rect 2486 430 2492 606
rect 2690 430 2700 610
rect 2760 430 2770 610
rect 2820 606 3140 656
rect 2820 430 2832 606
rect 2866 430 3090 606
rect 3124 430 3140 606
rect 1980 420 1990 430
rect 1944 418 1990 420
rect 2066 418 2112 430
rect 2324 418 2370 430
rect 2446 418 2492 430
rect 2704 418 2750 430
rect 1580 410 1720 418
rect 160 346 234 380
rect 402 346 480 380
rect 160 240 480 346
rect 602 380 794 386
rect 602 346 614 380
rect 782 346 794 380
rect 602 340 794 346
rect 982 380 1174 386
rect 982 346 994 380
rect 1162 346 1174 380
rect 982 340 1174 346
rect 1362 380 1554 386
rect 1362 346 1374 380
rect 1542 346 1554 380
rect 1362 340 1554 346
rect 1742 380 1934 386
rect 1742 346 1754 380
rect 1922 346 1934 380
rect 1742 340 1934 346
rect 2122 380 2314 386
rect 2122 346 2134 380
rect 2302 346 2314 380
rect 2122 340 2314 346
rect 2502 380 2694 386
rect 2502 346 2514 380
rect 2682 346 2694 380
rect 2502 340 2694 346
rect 2820 380 3140 430
rect 2820 346 2894 380
rect 3062 346 3140 380
rect 160 200 220 240
rect 440 210 480 240
rect 1088 240 1332 246
rect 1088 210 1100 240
rect 440 200 1100 210
rect 1320 210 1332 240
rect 2008 240 2252 246
rect 2008 210 2020 240
rect 1320 200 1580 210
rect 160 190 1580 200
rect 160 160 840 190
rect 160 40 200 160
rect 480 90 840 160
rect 940 90 1580 190
rect 480 70 1580 90
rect 1700 200 2020 210
rect 2240 210 2252 240
rect 2820 240 3140 346
rect 2820 210 2860 240
rect 2240 200 2340 210
rect 1700 70 2340 200
rect 2480 200 2860 210
rect 3080 200 3140 240
rect 2480 70 3140 200
rect 15720 160 15920 200
rect 480 40 3140 70
rect 160 0 3140 40
rect 14580 20 14600 160
rect 14700 140 17420 160
rect 14700 20 15640 140
rect 15900 20 17320 140
rect 17420 20 17430 140
rect 14580 0 17420 20
rect 16030 -20 16190 0
rect 60 -840 16100 -820
rect 60 -980 200 -840
rect -60 -1140 200 -980
rect 460 -860 16100 -840
rect 460 -880 15680 -860
rect 460 -920 5660 -880
rect 460 -1140 1060 -920
rect -60 -1180 1060 -1140
rect 60 -1200 1060 -1180
rect 1220 -1180 5660 -920
rect 5820 -1100 15680 -880
rect 15880 -1100 16100 -860
rect 5820 -1180 16100 -1100
rect 1220 -1200 16100 -1180
rect 60 -1260 16100 -1200
rect 4680 -1400 4880 -1380
rect 4680 -1500 4700 -1400
rect 4860 -1500 4880 -1400
rect 4680 -1800 4880 -1500
rect 13080 -1400 13280 -1380
rect 13080 -1500 13100 -1400
rect 13260 -1500 13280 -1400
rect 13080 -1800 13280 -1500
rect 14300 -1400 14500 -1380
rect 14300 -1500 14320 -1400
rect 14480 -1500 14500 -1400
rect 14300 -1600 14500 -1500
rect 14280 -1800 14480 -1600
<< via1 >>
rect 6940 33500 7260 33780
rect 5860 32440 6460 33060
rect 5840 31232 6440 31400
rect 5840 30835 6142 31232
rect 6142 30835 6180 31232
rect 6180 30835 6440 31232
rect 5840 30800 6440 30835
rect 1580 11320 1760 11460
rect 220 10660 500 10980
rect 1560 6560 1760 6760
rect 12880 6560 13080 6760
rect 1040 6400 1220 6560
rect 6300 6280 6460 6420
rect 6060 6180 6120 6260
rect 6580 6180 6640 6260
rect 7080 6180 7140 6260
rect 7460 6200 7520 6260
rect 8100 6180 8160 6260
rect 8620 6180 8680 6260
rect 9120 6180 9180 6260
rect 9520 6180 9580 6260
rect 10020 6180 10080 6260
rect 10540 6180 10600 6260
rect 10680 6180 10740 6260
rect 11320 6180 11380 6260
rect 11840 6180 11900 6260
rect 12360 6180 12420 6260
rect 6060 5988 6120 6000
rect 6060 5812 6066 5988
rect 6066 5812 6100 5988
rect 6100 5812 6120 5988
rect 6060 5800 6120 5812
rect 6300 5988 6360 6000
rect 6300 5812 6324 5988
rect 6324 5812 6358 5988
rect 6358 5812 6360 5988
rect 6300 5800 6360 5812
rect 6580 5988 6640 6000
rect 6580 5812 6582 5988
rect 6582 5812 6616 5988
rect 6616 5812 6640 5988
rect 6580 5800 6640 5812
rect 6820 5988 6880 6000
rect 6820 5812 6840 5988
rect 6840 5812 6874 5988
rect 6874 5812 6880 5988
rect 6820 5800 6880 5812
rect 7080 5988 7140 6000
rect 7080 5812 7098 5988
rect 7098 5812 7132 5988
rect 7132 5812 7140 5988
rect 7080 5800 7140 5812
rect 7340 5988 7400 6000
rect 7340 5812 7356 5988
rect 7356 5812 7390 5988
rect 7390 5812 7400 5988
rect 7340 5800 7400 5812
rect 7460 5988 7520 6000
rect 7460 5812 7468 5988
rect 7468 5812 7502 5988
rect 7502 5812 7520 5988
rect 7460 5800 7520 5812
rect 7700 5988 7760 6000
rect 7700 5812 7726 5988
rect 7726 5812 7760 5988
rect 7700 5800 7760 5812
rect 7840 5988 7900 6000
rect 7840 5812 7848 5988
rect 7848 5812 7882 5988
rect 7882 5812 7900 5988
rect 7840 5800 7900 5812
rect 8100 5988 8160 6000
rect 8100 5812 8106 5988
rect 8106 5812 8140 5988
rect 8140 5812 8160 5988
rect 8100 5800 8160 5812
rect 8360 5988 8420 6000
rect 8360 5812 8364 5988
rect 8364 5812 8398 5988
rect 8398 5812 8420 5988
rect 8360 5800 8420 5812
rect 8600 5988 8660 6000
rect 8600 5812 8622 5988
rect 8622 5812 8656 5988
rect 8656 5812 8660 5988
rect 8600 5800 8660 5812
rect 8860 5988 8920 6000
rect 8860 5812 8880 5988
rect 8880 5812 8914 5988
rect 8914 5812 8920 5988
rect 8860 5800 8920 5812
rect 9120 5988 9180 6000
rect 9120 5812 9138 5988
rect 9138 5812 9172 5988
rect 9172 5812 9180 5988
rect 9120 5800 9180 5812
rect 9260 5988 9320 6000
rect 9260 5812 9268 5988
rect 9268 5812 9302 5988
rect 9302 5812 9320 5988
rect 9260 5800 9320 5812
rect 9520 5988 9580 6000
rect 9520 5812 9526 5988
rect 9526 5812 9560 5988
rect 9560 5812 9580 5988
rect 9520 5800 9580 5812
rect 9780 5988 9840 6000
rect 9780 5812 9784 5988
rect 9784 5812 9818 5988
rect 9818 5812 9840 5988
rect 9780 5800 9840 5812
rect 10020 5988 10080 6000
rect 10020 5812 10042 5988
rect 10042 5812 10076 5988
rect 10076 5812 10080 5988
rect 10020 5800 10080 5812
rect 10280 5988 10340 6000
rect 10280 5812 10300 5988
rect 10300 5812 10334 5988
rect 10334 5812 10340 5988
rect 10280 5800 10340 5812
rect 10540 5988 10600 6000
rect 10540 5812 10558 5988
rect 10558 5812 10592 5988
rect 10592 5812 10600 5988
rect 10540 5800 10600 5812
rect 10680 5988 10740 6000
rect 10680 5812 10688 5988
rect 10688 5812 10722 5988
rect 10722 5812 10740 5988
rect 10680 5800 10740 5812
rect 11060 5988 11120 6000
rect 11060 5812 11068 5988
rect 11068 5812 11102 5988
rect 11102 5812 11120 5988
rect 11060 5800 11120 5812
rect 11320 5988 11380 6000
rect 11320 5812 11326 5988
rect 11326 5812 11360 5988
rect 11360 5812 11380 5988
rect 11320 5800 11380 5812
rect 11560 5988 11620 6000
rect 11560 5812 11584 5988
rect 11584 5812 11618 5988
rect 11618 5812 11620 5988
rect 11560 5800 11620 5812
rect 11840 5988 11900 6000
rect 11840 5812 11842 5988
rect 11842 5812 11876 5988
rect 11876 5812 11900 5988
rect 11840 5800 11900 5812
rect 12100 5988 12160 6000
rect 12100 5812 12134 5988
rect 12134 5812 12160 5988
rect 12100 5800 12160 5812
rect 12360 5988 12420 6000
rect 12360 5812 12392 5988
rect 12392 5812 12420 5988
rect 12360 5800 12420 5812
rect 10720 5719 10750 5740
rect 10750 5719 10780 5740
rect 10720 5680 10780 5719
rect 6300 5540 6360 5620
rect 6820 5540 6880 5620
rect 7220 5540 7280 5600
rect 7340 5540 7400 5620
rect 7840 5540 7900 5620
rect 8360 5540 8420 5620
rect 8860 5540 8920 5620
rect 9240 5540 9300 5620
rect 9760 5540 9820 5620
rect 10280 5540 10340 5620
rect 10600 5540 10660 5600
rect 11060 5540 11120 5620
rect 11560 5540 11620 5620
rect 12100 5540 12160 5620
rect 320 5300 400 5400
rect 1600 5300 1720 5400
rect 3500 5320 4000 5480
rect 4040 5300 4140 5400
rect 4380 5340 4560 5520
rect 6180 5420 6240 5480
rect 6340 5320 6400 5380
rect 6700 5320 6760 5380
rect 6860 5320 6920 5380
rect 7360 5320 7420 5380
rect 7880 5320 7940 5380
rect 8400 5320 8460 5380
rect 8920 5320 8980 5380
rect 9420 5320 9480 5380
rect 9940 5320 10000 5380
rect 10460 5320 10520 5380
rect 10980 5320 11040 5380
rect 11120 5340 11180 5400
rect 11600 5320 11660 5400
rect 6060 5200 6120 5260
rect 7100 5200 7160 5260
rect 7700 5200 7760 5260
rect 8140 5200 8200 5260
rect 9160 5200 9220 5260
rect 10200 5200 10260 5260
rect 11240 5200 11300 5260
rect 14300 5240 14440 5400
rect 17320 5700 17500 5880
rect 17360 5440 17460 5520
rect 11120 5120 11180 5160
rect 11120 5100 11180 5120
rect 6060 5070 6120 5080
rect 1600 4840 1720 4960
rect 2360 4592 2406 4800
rect 2406 4592 2440 4800
rect 2360 4580 2440 4592
rect 3280 4620 3380 4740
rect 4040 4840 4140 4960
rect 6060 4894 6096 5070
rect 6096 4894 6120 5070
rect 6060 4880 6120 4894
rect 6340 5070 6400 5080
rect 6340 4894 6354 5070
rect 6354 4894 6388 5070
rect 6388 4894 6400 5070
rect 6340 4880 6400 4894
rect 6580 5070 6640 5080
rect 6580 4894 6612 5070
rect 6612 4894 6640 5070
rect 6580 4880 6640 4894
rect 6860 5070 6920 5080
rect 6860 4894 6870 5070
rect 6870 4894 6904 5070
rect 6904 4894 6920 5070
rect 6860 4880 6920 4894
rect 7100 5070 7160 5080
rect 7100 4894 7128 5070
rect 7128 4894 7160 5070
rect 7100 4880 7160 4894
rect 7360 5070 7420 5080
rect 7360 4894 7386 5070
rect 7386 4894 7420 5070
rect 7360 4880 7420 4894
rect 7620 5070 7680 5080
rect 7620 4894 7644 5070
rect 7644 4894 7678 5070
rect 7678 4894 7680 5070
rect 7620 4880 7680 4894
rect 7880 5070 7940 5080
rect 7880 4894 7902 5070
rect 7902 4894 7936 5070
rect 7936 4894 7940 5070
rect 7880 4880 7940 4894
rect 8140 5070 8200 5080
rect 8140 4894 8160 5070
rect 8160 4894 8194 5070
rect 8194 4894 8200 5070
rect 8140 4880 8200 4894
rect 8400 5070 8460 5080
rect 8400 4894 8418 5070
rect 8418 4894 8452 5070
rect 8452 4894 8460 5070
rect 8400 4880 8460 4894
rect 8660 4894 8676 5070
rect 8676 4894 8710 5070
rect 8710 4894 8720 5070
rect 8660 4890 8720 4894
rect 8920 5070 8980 5080
rect 8920 4894 8934 5070
rect 8934 4894 8968 5070
rect 8968 4894 8980 5070
rect 8920 4880 8980 4894
rect 9160 5070 9220 5080
rect 9160 4894 9192 5070
rect 9192 4894 9220 5070
rect 9160 4880 9220 4894
rect 9420 5070 9480 5080
rect 9420 4894 9450 5070
rect 9450 4894 9480 5070
rect 9420 4880 9480 4894
rect 9680 5070 9740 5080
rect 9680 4894 9708 5070
rect 9708 4894 9740 5070
rect 9680 4880 9740 4894
rect 9940 5070 10000 5080
rect 9940 4894 9966 5070
rect 9966 4894 10000 5070
rect 9940 4880 10000 4894
rect 10200 5070 10260 5080
rect 10200 4894 10224 5070
rect 10224 4894 10258 5070
rect 10258 4894 10260 5070
rect 10200 4880 10260 4894
rect 10460 5070 10520 5080
rect 10460 4894 10482 5070
rect 10482 4894 10516 5070
rect 10516 4894 10520 5070
rect 10460 4880 10520 4894
rect 10720 4894 10740 5070
rect 10740 4894 10774 5070
rect 10774 4894 10780 5070
rect 10720 4880 10780 4894
rect 10980 4894 10998 5060
rect 10998 4894 11032 5060
rect 11032 4894 11040 5060
rect 10980 4880 11040 4894
rect 11240 4894 11256 5060
rect 11256 4894 11290 5060
rect 11290 4894 11300 5060
rect 11240 4880 11300 4894
rect 6180 4800 6240 4860
rect 6580 4700 6640 4760
rect 7620 4700 7680 4760
rect 8660 4700 8720 4760
rect 9680 4700 9740 4760
rect 10720 4700 10780 4760
rect 2620 4533 2720 4540
rect 2620 4499 2720 4533
rect 2620 4480 2720 4499
rect 4700 4480 4880 4640
rect 6180 4540 6240 4600
rect 6820 4500 6880 4560
rect 7220 4500 7280 4560
rect 7880 4500 7940 4560
rect 8900 4500 8960 4560
rect 9940 4500 10000 4560
rect 10960 4500 11020 4560
rect 12000 4500 12060 4560
rect 7360 4380 7420 4440
rect 8400 4380 8460 4440
rect 9420 4380 9480 4440
rect 10440 4380 10500 4440
rect 10600 4380 10660 4440
rect 11480 4380 11540 4440
rect 11600 4380 11660 4440
rect 320 4271 400 4300
rect 320 4220 388 4271
rect 388 4220 400 4271
rect 2360 4200 2440 4300
rect 2920 4180 3020 4280
rect 6180 4236 6240 4240
rect 6180 4060 6190 4236
rect 6190 4060 6224 4236
rect 6224 4060 6240 4236
rect 6440 4060 6448 4200
rect 6448 4060 6482 4200
rect 6482 4060 6500 4200
rect 6700 4060 6706 4200
rect 6706 4060 6740 4200
rect 6740 4060 6760 4200
rect 6840 4060 6852 4220
rect 6852 4060 6886 4220
rect 6886 4060 6900 4220
rect 7100 4060 7110 4220
rect 7110 4060 7144 4220
rect 7144 4060 7160 4220
rect 7360 4060 7368 4220
rect 7368 4060 7402 4220
rect 7402 4060 7420 4220
rect 7620 4060 7626 4220
rect 7626 4060 7660 4220
rect 7660 4060 7680 4220
rect 7880 4060 7884 4220
rect 7884 4060 7918 4220
rect 7918 4060 7940 4220
rect 8140 4060 8142 4220
rect 8142 4060 8176 4220
rect 8176 4060 8200 4220
rect 8400 4060 8434 4220
rect 8434 4060 8460 4220
rect 8640 4060 8658 4220
rect 8658 4060 8692 4220
rect 8692 4060 8700 4220
rect 8900 4060 8916 4220
rect 8916 4060 8950 4220
rect 8950 4060 8960 4220
rect 9160 4060 9174 4220
rect 9174 4060 9208 4220
rect 9208 4060 9220 4220
rect 9420 4060 9432 4220
rect 9432 4060 9466 4220
rect 9466 4060 9480 4220
rect 9680 4060 9690 4220
rect 9690 4060 9724 4220
rect 9724 4060 9740 4220
rect 9940 4060 9948 4220
rect 9948 4060 9982 4220
rect 9982 4060 10000 4220
rect 10200 4060 10206 4220
rect 10206 4060 10240 4220
rect 10240 4060 10260 4220
rect 10440 4060 10464 4220
rect 10464 4060 10498 4220
rect 10498 4060 10500 4220
rect 10700 4060 10722 4220
rect 10722 4060 10756 4220
rect 10756 4060 10760 4220
rect 10960 4060 10980 4220
rect 10980 4060 11014 4220
rect 11014 4060 11020 4220
rect 11220 4060 11238 4220
rect 11238 4060 11272 4220
rect 11272 4060 11280 4220
rect 11480 4060 11496 4220
rect 11496 4060 11530 4220
rect 11530 4060 11540 4220
rect 11740 4060 11754 4220
rect 11754 4060 11788 4220
rect 11788 4060 11800 4220
rect 12000 4060 12012 4220
rect 12012 4060 12046 4220
rect 12046 4060 12060 4220
rect 14320 4160 14460 4320
rect 15860 4020 15940 4380
rect 840 3853 940 3860
rect 840 3819 940 3853
rect 840 3800 940 3819
rect 2620 3853 2720 3860
rect 2620 3819 2630 3853
rect 2630 3819 2720 3853
rect 2620 3800 2720 3819
rect 5660 3700 5840 3900
rect 6440 3840 6500 3900
rect 7100 3840 7160 3900
rect 7620 3840 7680 3900
rect 8140 3840 8200 3900
rect 8640 3840 8700 3900
rect 9160 3840 9220 3900
rect 9680 3840 9740 3900
rect 10200 3840 10260 3900
rect 10700 3840 10760 3900
rect 11220 3840 11280 3900
rect 11740 3840 11800 3900
rect 16780 3880 16860 3940
rect 15860 3720 15940 3800
rect 17180 3720 17260 3820
rect 2620 3420 2720 3540
rect 17180 3494 17240 3520
rect 17180 3460 17208 3494
rect 17208 3460 17240 3494
rect 12880 3240 13080 3440
rect 16900 3260 16970 3370
rect 2620 2613 2700 2780
rect 3280 2940 3360 3040
rect 3360 2940 3400 3040
rect 4380 2900 4560 3100
rect 14340 2960 14460 3080
rect 14340 2940 14430 2960
rect 14430 2940 14460 2960
rect 17080 2840 17140 3420
rect 17360 3300 17400 3380
rect 17400 3300 17440 3380
rect 17360 3180 17400 3260
rect 17400 3180 17440 3260
rect 17360 3040 17400 3120
rect 17400 3040 17440 3120
rect 17360 2900 17400 2980
rect 17400 2900 17440 2980
rect 2620 2580 2700 2613
rect 13080 2580 13260 2760
rect 14890 2650 14970 2660
rect 14890 2610 14900 2650
rect 14900 2610 14960 2650
rect 14960 2610 14970 2650
rect 14890 2590 14970 2610
rect 15340 2655 15400 2660
rect 15340 2621 15359 2655
rect 15359 2621 15393 2655
rect 15393 2621 15400 2655
rect 16900 2660 16980 2740
rect 17200 2732 17208 2760
rect 17208 2732 17242 2760
rect 17242 2732 17260 2760
rect 17200 2700 17260 2732
rect 15340 2600 15400 2621
rect 16780 2560 16860 2620
rect 2040 2420 2100 2480
rect 2920 2420 3020 2480
rect 14620 2485 14700 2500
rect 14620 2451 14627 2485
rect 14627 2451 14661 2485
rect 14661 2451 14700 2485
rect 14620 2420 14700 2451
rect 17200 2406 17260 2440
rect 17200 2380 17208 2406
rect 17208 2380 17242 2406
rect 17242 2380 17260 2406
rect 540 2240 600 2320
rect 840 2240 940 2300
rect 1180 2240 1240 2320
rect 1300 2280 1360 2360
rect 1940 2280 2000 2360
rect 2620 2280 2720 2360
rect 14900 2320 14960 2380
rect 17060 2310 17120 2370
rect 2700 2080 2760 2160
rect 2920 2080 3000 2160
rect 14340 2020 14460 2200
rect 15340 2100 15400 2160
rect 17320 2140 17360 2280
rect 17360 2140 17400 2280
rect 17400 2140 17420 2280
rect 2680 1944 2760 1980
rect 2680 1920 2682 1944
rect 2682 1920 2760 1944
rect 540 1860 600 1870
rect 540 1690 552 1860
rect 552 1690 586 1860
rect 586 1690 600 1860
rect 820 1860 960 1870
rect 820 1684 844 1860
rect 844 1684 932 1860
rect 932 1684 960 1860
rect 1180 1860 1240 1870
rect 1180 1690 1190 1860
rect 1190 1690 1224 1860
rect 1224 1690 1240 1860
rect 1300 1690 1312 1850
rect 1312 1690 1346 1850
rect 1346 1690 1360 1850
rect 820 1670 960 1684
rect 1580 1690 1604 1830
rect 1604 1690 1680 1830
rect 1920 1684 1950 1860
rect 1950 1684 1980 1860
rect 1920 1680 1980 1684
rect 2040 1860 2120 1870
rect 2040 1684 2072 1860
rect 2072 1684 2106 1860
rect 2106 1684 2120 1860
rect 2040 1670 2120 1684
rect 2340 1690 2364 1850
rect 2364 1690 2452 1850
rect 2452 1690 2460 1850
rect 2680 1684 2710 1850
rect 2710 1684 2740 1850
rect 2680 1670 2740 1684
rect 540 1442 600 1450
rect 540 1266 552 1442
rect 552 1266 586 1442
rect 586 1266 600 1442
rect 540 1250 600 1266
rect 820 1442 960 1450
rect 820 1266 844 1442
rect 844 1266 932 1442
rect 932 1266 960 1442
rect 1180 1442 1240 1450
rect 1180 1270 1190 1442
rect 1190 1270 1224 1442
rect 1224 1270 1240 1442
rect 1300 1270 1312 1430
rect 1312 1270 1346 1430
rect 1346 1270 1360 1430
rect 820 1250 960 1266
rect 1600 1270 1604 1410
rect 1604 1270 1692 1410
rect 1692 1270 1700 1410
rect 1920 1266 1950 1440
rect 1950 1266 1980 1440
rect 1920 1260 1980 1266
rect 2060 1442 2140 1450
rect 2060 1266 2072 1442
rect 2072 1266 2106 1442
rect 2106 1266 2140 1442
rect 2060 1250 2140 1266
rect 2340 1270 2364 1430
rect 2364 1270 2452 1430
rect 2452 1270 2460 1430
rect 2700 1442 2760 1450
rect 2700 1270 2710 1442
rect 2710 1270 2744 1442
rect 2744 1270 2760 1442
rect 540 1024 600 1030
rect 540 850 552 1024
rect 552 850 586 1024
rect 586 850 600 1024
rect 820 1024 960 1030
rect 820 848 844 1024
rect 844 848 932 1024
rect 932 848 960 1024
rect 1180 1024 1240 1030
rect 1180 850 1190 1024
rect 1190 850 1224 1024
rect 1224 850 1240 1024
rect 1300 850 1312 1010
rect 1312 850 1346 1010
rect 1346 850 1360 1010
rect 820 830 960 848
rect 1600 850 1604 990
rect 1604 850 1692 990
rect 1692 850 1700 990
rect 1920 848 1950 1020
rect 1950 848 1980 1020
rect 2060 1024 2120 1030
rect 2060 850 2072 1024
rect 2072 850 2106 1024
rect 2106 850 2120 1024
rect 1920 840 1980 848
rect 2340 850 2364 1010
rect 2364 850 2452 1010
rect 2452 850 2460 1010
rect 2700 1024 2760 1030
rect 2700 850 2710 1024
rect 2710 850 2744 1024
rect 2744 850 2760 1024
rect 540 606 600 610
rect 540 430 552 606
rect 552 430 586 606
rect 586 430 600 606
rect 820 606 960 610
rect 820 430 844 606
rect 844 430 932 606
rect 932 430 960 606
rect 1180 606 1240 610
rect 1180 430 1190 606
rect 1190 430 1224 606
rect 1224 430 1240 606
rect 1300 430 1312 590
rect 1312 430 1346 590
rect 1346 430 1360 590
rect 1600 430 1604 570
rect 1604 430 1692 570
rect 1692 430 1700 570
rect 1920 430 1950 600
rect 1950 430 1980 600
rect 2060 606 2120 610
rect 2060 430 2072 606
rect 2072 430 2106 606
rect 2106 430 2120 606
rect 2340 430 2364 590
rect 2364 430 2452 590
rect 2452 430 2460 590
rect 2700 606 2760 610
rect 2700 430 2710 606
rect 2710 430 2744 606
rect 2744 430 2760 606
rect 1920 420 1980 430
rect 200 40 480 160
rect 840 90 940 190
rect 1580 70 1700 210
rect 2340 70 2480 210
rect 14600 20 14700 160
rect 15640 20 15900 140
rect 17320 20 17420 140
rect 200 -1140 460 -840
rect 1060 -1200 1220 -920
rect 5660 -1180 5820 -880
rect 15680 -1100 15880 -860
rect 4700 -1500 4860 -1400
rect 13100 -1500 13260 -1400
rect 14320 -1500 14480 -1400
<< metal2 >>
rect 6940 33780 7260 33790
rect 6940 33490 7260 33500
rect 5860 33060 6460 33070
rect 5860 32430 6460 32440
rect 5840 31400 6440 31410
rect 5840 30790 6440 30800
rect 1560 11460 1780 11500
rect 1560 11320 1580 11460
rect 1760 11320 1780 11460
rect 220 10980 500 10990
rect 220 10650 500 10660
rect 1560 6760 1780 11320
rect 1040 6560 1220 6570
rect 1760 6560 1780 6760
rect 12880 6760 13100 6780
rect 13080 6560 13100 6760
rect 1560 6550 1760 6560
rect 1040 6390 1220 6400
rect 6300 6420 6460 6430
rect 6300 6270 6460 6280
rect 6060 6260 6120 6270
rect 6060 6000 6120 6180
rect 6580 6260 6640 6270
rect 6060 5790 6120 5800
rect 6300 6000 6360 6010
rect 6300 5620 6360 5800
rect 6580 6000 6640 6180
rect 7080 6260 7140 6270
rect 6580 5790 6640 5800
rect 6820 6000 6880 6010
rect 4360 5520 4560 5540
rect 6300 5530 6360 5540
rect 6820 5620 6880 5800
rect 7080 6000 7140 6180
rect 7460 6260 7520 6270
rect 7080 5790 7140 5800
rect 7340 6000 7400 6010
rect 7340 5620 7400 5800
rect 7460 6000 7520 6200
rect 8100 6260 8160 6270
rect 7460 5790 7520 5800
rect 7700 6000 7760 6010
rect 6820 5530 6880 5540
rect 7220 5600 7280 5620
rect 3500 5480 4000 5490
rect 320 5400 400 5410
rect 320 4300 400 5300
rect 1600 5400 1720 5410
rect 3500 5310 4000 5320
rect 4040 5400 4140 5410
rect 1600 4960 1720 5300
rect 1600 4830 1720 4840
rect 4040 4960 4140 5300
rect 4040 4830 4140 4840
rect 4360 5340 4380 5520
rect 320 4210 400 4220
rect 2360 4800 2440 4810
rect 2360 4300 2440 4580
rect 3280 4740 3400 4760
rect 3380 4620 3400 4740
rect 2360 4190 2440 4200
rect 2620 4540 2720 4550
rect 840 3860 940 3870
rect 540 2320 600 2330
rect 540 1870 600 2240
rect 840 2300 940 3800
rect 2620 3860 2720 4480
rect 2620 3540 2720 3800
rect 2620 2780 2720 3420
rect 2700 2580 2720 2780
rect 2040 2480 2100 2490
rect 1300 2360 1360 2370
rect 840 2230 940 2240
rect 1180 2320 1240 2330
rect 540 1450 600 1690
rect 540 1030 600 1250
rect 540 610 600 850
rect 540 410 600 430
rect 820 1870 960 1880
rect 820 1450 960 1670
rect 820 1030 960 1250
rect 820 610 960 830
rect 820 190 960 430
rect 1180 1870 1240 2240
rect 1180 1450 1240 1690
rect 1180 1030 1240 1270
rect 1180 610 1240 850
rect 1180 410 1240 430
rect 1300 1850 1360 2280
rect 1940 2360 2000 2370
rect 1940 1870 2000 2280
rect 1920 1860 2000 1870
rect 1300 1430 1360 1690
rect 1300 1010 1360 1270
rect 1300 590 1360 850
rect 1300 410 1360 430
rect 1580 1830 1700 1850
rect 1680 1690 1700 1830
rect 1580 1410 1700 1690
rect 1980 1680 2000 1860
rect 1920 1670 2000 1680
rect 1940 1450 2000 1670
rect 1580 1270 1600 1410
rect 1580 990 1700 1270
rect 1920 1440 2000 1450
rect 1980 1260 2000 1440
rect 1920 1250 2000 1260
rect 1940 1030 2000 1250
rect 1580 850 1600 990
rect 1580 570 1700 850
rect 1920 1020 2000 1030
rect 1980 840 2000 1020
rect 1920 830 2000 840
rect 1940 610 2000 830
rect 1580 430 1600 570
rect 160 160 500 180
rect 160 40 200 160
rect 480 40 500 160
rect 820 90 840 190
rect 940 90 960 190
rect 820 70 960 90
rect 1580 210 1700 430
rect 1920 600 2000 610
rect 1980 420 2000 600
rect 1920 410 2000 420
rect 2040 1880 2100 2420
rect 2620 2360 2720 2580
rect 2620 2270 2720 2280
rect 2920 4280 3020 4290
rect 2920 2480 3020 4180
rect 3280 3040 3400 4620
rect 3280 2930 3400 2940
rect 4360 3100 4560 5340
rect 6180 5480 6240 5490
rect 6060 5260 6120 5280
rect 6060 5080 6120 5200
rect 6060 4870 6120 4880
rect 6180 4860 6240 5420
rect 6340 5380 6400 5390
rect 6340 5080 6400 5320
rect 6700 5380 6760 5390
rect 6340 4870 6400 4880
rect 6580 5080 6640 5090
rect 6180 4790 6240 4800
rect 6580 4760 6640 4880
rect 6580 4690 6640 4700
rect 4360 2900 4380 3100
rect 4380 2890 4560 2900
rect 4660 4640 4880 4680
rect 4660 4480 4700 4640
rect 2920 2390 3020 2420
rect 2700 2160 2760 2170
rect 2700 1990 2760 2080
rect 2920 2160 3000 2390
rect 2920 2070 3000 2080
rect 2680 1980 2760 1990
rect 2680 1910 2760 1920
rect 2040 1870 2120 1880
rect 2040 1660 2120 1670
rect 2340 1850 2480 1870
rect 2700 1860 2760 1910
rect 2460 1690 2480 1850
rect 2040 1460 2100 1660
rect 2040 1450 2140 1460
rect 2040 1250 2060 1450
rect 2040 1240 2140 1250
rect 2340 1430 2480 1690
rect 2680 1850 2760 1860
rect 2740 1670 2760 1850
rect 2680 1660 2760 1670
rect 2460 1270 2480 1430
rect 2040 1040 2100 1240
rect 2040 1030 2120 1040
rect 2040 850 2060 1030
rect 2040 840 2120 850
rect 2340 1010 2480 1270
rect 2460 850 2480 1010
rect 2040 620 2100 840
rect 2040 610 2120 620
rect 2040 430 2060 610
rect 2040 420 2120 430
rect 2340 590 2480 850
rect 2460 430 2480 590
rect 2040 350 2100 420
rect 1580 60 1700 70
rect 2340 210 2480 430
rect 2700 1450 2760 1660
rect 2700 1030 2760 1270
rect 2700 610 2760 850
rect 2700 370 2760 430
rect 2340 60 2480 70
rect 160 -840 500 40
rect 160 -1140 200 -840
rect 460 -1140 500 -840
rect 160 -1180 500 -1140
rect 1060 -920 1220 -910
rect 1060 -1210 1220 -1200
rect 4660 -1400 4880 4480
rect 6180 4600 6240 4610
rect 6180 4240 6240 4540
rect 6180 4050 6240 4060
rect 6440 4200 6500 4210
rect 5640 3900 5840 3920
rect 5640 3700 5660 3900
rect 6440 3900 6500 4060
rect 6700 4200 6760 5320
rect 6860 5380 6920 5390
rect 6860 5080 6920 5320
rect 6860 4870 6920 4880
rect 7100 5260 7160 5270
rect 7100 5080 7160 5200
rect 7100 4870 7160 4880
rect 6700 4050 6760 4060
rect 6820 4560 6880 4570
rect 6820 4230 6880 4500
rect 7220 4560 7280 5540
rect 7340 5530 7400 5540
rect 7360 5380 7420 5390
rect 7360 5080 7420 5320
rect 7700 5260 7760 5800
rect 7840 6000 7900 6010
rect 7840 5620 7900 5800
rect 8100 6000 8160 6180
rect 8620 6260 8680 6270
rect 8620 6010 8680 6180
rect 9120 6260 9180 6270
rect 8100 5790 8160 5800
rect 8360 6000 8420 6010
rect 7840 5530 7900 5540
rect 8360 5620 8420 5800
rect 8600 6000 8680 6010
rect 8660 5800 8680 6000
rect 8860 6000 8920 6010
rect 8600 5790 8660 5800
rect 8360 5530 8420 5540
rect 8860 5620 8920 5800
rect 9120 6000 9180 6180
rect 9520 6260 9580 6270
rect 9260 6000 9320 6010
rect 9120 5790 9180 5800
rect 9240 5800 9260 6000
rect 9240 5790 9320 5800
rect 9520 6000 9580 6180
rect 10020 6260 10080 6270
rect 9780 6000 9840 6010
rect 9520 5790 9580 5800
rect 9760 5800 9780 6000
rect 9760 5790 9840 5800
rect 10020 6000 10080 6180
rect 10540 6260 10600 6270
rect 10020 5790 10080 5800
rect 10280 6000 10340 6010
rect 8860 5530 8920 5540
rect 9240 5620 9300 5790
rect 9240 5530 9300 5540
rect 9760 5620 9820 5790
rect 9760 5530 9820 5540
rect 10280 5620 10340 5800
rect 10540 6000 10600 6180
rect 10540 5790 10600 5800
rect 10680 6260 10740 6270
rect 10680 6000 10740 6180
rect 11320 6260 11380 6270
rect 10680 5790 10740 5800
rect 11060 6000 11120 6010
rect 10720 5740 10780 5760
rect 10280 5520 10340 5540
rect 10600 5600 10660 5610
rect 7700 5190 7760 5200
rect 7880 5380 7940 5390
rect 7360 4870 7420 4880
rect 7620 5080 7680 5090
rect 7620 4760 7680 4880
rect 7880 5080 7940 5320
rect 8400 5380 8460 5390
rect 7880 4870 7940 4880
rect 8140 5260 8200 5270
rect 8140 5080 8200 5200
rect 8140 4870 8200 4880
rect 8400 5080 8460 5320
rect 8920 5380 8980 5390
rect 8920 5080 8980 5320
rect 9420 5380 9480 5390
rect 8400 4870 8460 4880
rect 8660 5070 8720 5080
rect 7620 4690 7680 4700
rect 8660 4760 8720 4890
rect 8920 4870 8980 4880
rect 9160 5260 9220 5270
rect 9160 5080 9220 5200
rect 9160 4870 9220 4880
rect 9420 5080 9480 5320
rect 9940 5380 10000 5390
rect 9420 4870 9480 4880
rect 9680 5080 9740 5090
rect 8660 4690 8720 4700
rect 9680 4760 9740 4880
rect 9940 5080 10000 5320
rect 10460 5380 10520 5390
rect 9940 4870 10000 4880
rect 10200 5260 10260 5270
rect 10200 5080 10260 5200
rect 10200 4870 10260 4880
rect 10460 5080 10520 5320
rect 10460 4870 10520 4880
rect 9680 4690 9740 4700
rect 7220 4490 7280 4500
rect 7880 4560 7940 4570
rect 7360 4440 7420 4450
rect 6820 4220 6900 4230
rect 6820 4060 6840 4220
rect 6820 4050 6900 4060
rect 7100 4220 7160 4230
rect 6440 3830 6500 3840
rect 5640 -880 5840 3700
rect 6820 3520 6880 4050
rect 7100 3900 7160 4060
rect 7360 4220 7420 4380
rect 7360 4050 7420 4060
rect 7620 4220 7680 4230
rect 7100 3830 7160 3840
rect 7620 3900 7680 4060
rect 7880 4220 7940 4500
rect 8900 4560 8960 4570
rect 8400 4440 8460 4450
rect 7880 4050 7940 4060
rect 8140 4220 8200 4230
rect 7620 3830 7680 3840
rect 8140 3900 8200 4060
rect 8400 4220 8460 4380
rect 8400 4050 8460 4060
rect 8640 4220 8700 4230
rect 8140 3830 8200 3840
rect 8640 3900 8700 4060
rect 8900 4220 8960 4500
rect 9940 4560 10000 4570
rect 9420 4440 9480 4450
rect 8900 4040 8960 4060
rect 9160 4220 9220 4230
rect 8640 3830 8700 3840
rect 9160 3900 9220 4060
rect 9420 4220 9480 4380
rect 9420 4040 9480 4060
rect 9680 4220 9740 4230
rect 9160 3830 9220 3840
rect 9680 3900 9740 4060
rect 9940 4220 10000 4500
rect 10440 4440 10500 4450
rect 9940 4040 10000 4060
rect 10200 4220 10260 4230
rect 9680 3830 9740 3840
rect 10200 3900 10260 4060
rect 10440 4220 10500 4380
rect 10600 4440 10660 5540
rect 10720 5080 10780 5680
rect 11060 5620 11120 5800
rect 11320 6000 11380 6180
rect 11840 6260 11900 6270
rect 11320 5790 11380 5800
rect 11560 6000 11620 6010
rect 11060 5530 11120 5540
rect 11560 5620 11620 5800
rect 11840 6000 11900 6180
rect 12360 6260 12420 6270
rect 11840 5790 11900 5800
rect 12100 6000 12160 6010
rect 11560 5530 11620 5540
rect 12100 5620 12160 5800
rect 12360 6000 12420 6180
rect 12360 5790 12420 5800
rect 12100 5530 12160 5540
rect 11120 5400 11180 5410
rect 10710 5070 10780 5080
rect 10710 4880 10720 5070
rect 10720 4760 10780 4880
rect 10980 5380 11040 5390
rect 10980 5060 11040 5320
rect 11120 5160 11180 5340
rect 11600 5400 11660 5410
rect 11120 5090 11180 5100
rect 11240 5260 11300 5270
rect 10980 4870 11040 4880
rect 11240 5060 11300 5200
rect 11240 4870 11300 4880
rect 10720 4690 10780 4700
rect 10600 4360 10660 4380
rect 10960 4560 11020 4570
rect 10440 4040 10500 4060
rect 10700 4220 10760 4230
rect 10200 3830 10260 3840
rect 10700 3900 10760 4060
rect 10960 4220 11020 4500
rect 11480 4440 11540 4450
rect 10960 4040 11020 4060
rect 11220 4220 11280 4230
rect 10700 3830 10760 3840
rect 11220 3900 11280 4060
rect 11480 4220 11540 4380
rect 11480 4040 11540 4060
rect 11600 4440 11660 5320
rect 11220 3830 11280 3840
rect 11600 3780 11660 4380
rect 12000 4560 12060 4570
rect 11740 4220 11800 4230
rect 11740 3900 11800 4060
rect 12000 4220 12060 4500
rect 12000 4040 12060 4060
rect 11740 3830 11800 3840
rect 11600 3690 11660 3700
rect 6820 3430 6880 3440
rect 12880 3440 13100 6560
rect 17320 5880 17500 5890
rect 17320 5690 17500 5700
rect 17360 5520 17460 5530
rect 17340 5440 17360 5520
rect 14280 5400 14460 5420
rect 14280 5240 14300 5400
rect 14440 5240 14460 5400
rect 14280 4320 14460 5240
rect 14280 4160 14320 4320
rect 14280 4140 14460 4160
rect 15860 4380 15960 4400
rect 15940 4020 15960 4380
rect 15860 3800 15960 4020
rect 15940 3720 15960 3800
rect 15860 3680 15960 3720
rect 16780 3940 16860 3950
rect 13080 3240 13100 3440
rect 12880 3230 13080 3240
rect 14300 3080 14500 3120
rect 14300 2940 14340 3080
rect 14460 2940 14500 3080
rect 5640 -1180 5660 -880
rect 5820 -1180 5840 -880
rect 5640 -1260 5840 -1180
rect 13080 2760 13280 2780
rect 13260 2580 13280 2760
rect 4660 -1500 4700 -1400
rect 4860 -1500 4880 -1400
rect 4660 -1520 4880 -1500
rect 13080 -1400 13280 2580
rect 13080 -1500 13100 -1400
rect 13260 -1500 13280 -1400
rect 13080 -1520 13280 -1500
rect 14300 2200 14500 2940
rect 14890 2660 14970 2670
rect 14890 2580 14970 2590
rect 15340 2660 15400 2670
rect 14620 2500 14700 2510
rect 14300 2020 14340 2200
rect 14460 2020 14500 2200
rect 14300 -1400 14500 2020
rect 14600 2420 14620 2500
rect 14600 160 14700 2420
rect 14900 2390 14940 2580
rect 14900 2380 14960 2390
rect 14900 2310 14960 2320
rect 15340 2160 15400 2600
rect 16780 2620 16860 3880
rect 17180 3820 17300 3830
rect 17180 3690 17300 3700
rect 17180 3520 17260 3690
rect 17240 3460 17260 3520
rect 17180 3450 17240 3460
rect 17080 3420 17140 3430
rect 16900 3370 16970 3380
rect 16900 2750 16970 3260
rect 17340 3380 17460 5440
rect 17340 3300 17360 3380
rect 17440 3300 17460 3380
rect 17340 3260 17460 3300
rect 17340 3180 17360 3260
rect 17440 3180 17460 3260
rect 17340 3120 17460 3180
rect 17340 3040 17360 3120
rect 17440 3040 17460 3120
rect 17340 2980 17460 3040
rect 17340 2900 17360 2980
rect 17440 2900 17460 2980
rect 17340 2840 17460 2900
rect 16900 2740 16980 2750
rect 16900 2650 16980 2660
rect 16780 2550 16860 2560
rect 17080 2380 17140 2840
rect 17060 2370 17140 2380
rect 17200 2760 17260 2770
rect 17200 2440 17260 2700
rect 17200 2370 17260 2380
rect 17120 2310 17140 2370
rect 17060 2300 17140 2310
rect 17080 2140 17140 2300
rect 17320 2280 17420 2300
rect 15340 2090 15400 2100
rect 14600 10 14700 20
rect 15600 140 15940 200
rect 15600 20 15640 140
rect 15900 20 15940 140
rect 15600 -860 15940 20
rect 17320 140 17420 2140
rect 17320 10 17420 20
rect 15600 -1100 15680 -860
rect 15880 -1100 15940 -860
rect 15600 -1180 15940 -1100
rect 14300 -1500 14320 -1400
rect 14480 -1500 14500 -1400
rect 14300 -1520 14500 -1500
<< via2 >>
rect 6940 33500 7260 33780
rect 5860 32440 6460 33060
rect 5840 30800 6440 31400
rect 220 10660 500 10980
rect 1040 6400 1220 6560
rect 6300 6280 6460 6420
rect 3500 5320 4000 5480
rect 1060 -1200 1220 -920
rect 11600 3700 11660 3780
rect 6820 3440 6880 3520
rect 17320 5700 17500 5880
rect 17180 3720 17260 3820
rect 17260 3720 17300 3820
rect 17180 3700 17300 3720
rect 17320 40 17420 140
<< metal3 >>
rect 6930 33780 7270 33785
rect 6930 33500 6940 33780
rect 7260 33500 7270 33780
rect 6930 33495 7270 33500
rect 5850 33060 6470 33065
rect 5850 32440 5860 33060
rect 6460 32440 6470 33060
rect 5850 32435 6470 32440
rect 5830 31400 6450 31405
rect 5830 30800 5840 31400
rect 6440 30800 6450 31400
rect 5830 30795 6450 30800
rect 210 10980 510 10985
rect 210 10660 220 10980
rect 500 10660 510 10980
rect 210 10655 510 10660
rect 120 9040 22338 9120
rect 120 6840 160 9040
rect 600 8900 22338 9040
rect 600 6880 20200 8900
rect 22120 6880 22338 8900
rect 600 6840 22338 6880
rect 120 6760 22338 6840
rect 1040 6565 1240 6580
rect 1030 6560 1240 6565
rect 1030 6400 1040 6560
rect 1220 6400 1240 6560
rect 6290 6420 6470 6425
rect 1030 6395 1240 6400
rect 1040 -920 1240 6395
rect 6260 6280 6300 6420
rect 6460 6400 7260 6420
rect 6460 6280 6900 6400
rect 7240 6280 7260 6400
rect 6290 6275 6470 6280
rect 6980 5920 17520 5940
rect 6980 5720 7000 5920
rect 7260 5880 17520 5920
rect 7260 5720 17320 5880
rect 6980 5700 17320 5720
rect 17500 5700 17520 5880
rect 17310 5695 17510 5700
rect 3490 5480 4010 5485
rect 3480 5320 3500 5480
rect 4000 5320 6920 5480
rect 3480 5300 6920 5320
rect 7240 5300 7250 5480
rect 3480 5280 7220 5300
rect 17160 3820 17320 3840
rect 11590 3780 11670 3785
rect 11590 3760 11600 3780
rect 11560 3700 11600 3760
rect 11660 3760 11670 3780
rect 11660 3740 12200 3760
rect 11660 3700 11960 3740
rect 11560 3680 11960 3700
rect 11950 3540 11960 3680
rect 12260 3540 12270 3740
rect 17160 3700 17180 3820
rect 17300 3700 17320 3820
rect 17160 3680 17320 3700
rect 6810 3520 6890 3525
rect 6010 3440 6020 3520
rect 6140 3440 6820 3520
rect 6880 3440 6890 3520
rect 6810 3435 6890 3440
rect 17300 140 17440 160
rect 17280 40 17320 140
rect 17420 40 17440 140
rect 17720 124 23240 5852
rect 17720 60 17748 124
rect 23212 60 23240 124
rect 17720 40 23240 60
rect 17280 20 17440 40
rect 1040 -1200 1060 -920
rect 1220 -1200 1240 -920
rect 1040 -1260 1240 -1200
<< via3 >>
rect 6940 33500 7260 33780
rect 5860 32440 6460 33060
rect 5840 30800 6440 31400
rect 220 10660 500 10980
rect 160 6840 600 9040
rect 20200 6880 22120 8900
rect 6900 6280 7240 6400
rect 7000 5720 7260 5920
rect 6920 5300 7240 5480
rect 11960 3540 12260 3740
rect 17180 3700 17300 3820
rect 6020 3440 6140 3520
rect 17320 40 17420 140
rect 17748 60 23212 124
<< mimcap >>
rect 17760 5772 23200 5812
rect 17760 412 17800 5772
rect 23160 412 23200 5772
rect 17760 372 23200 412
<< mimcapcontact >>
rect 17800 412 23160 5772
<< metal4 >>
rect 6900 33780 7280 33860
rect 6900 33500 6940 33780
rect 7260 33500 7280 33780
rect 5859 33060 6461 33061
rect 122 32999 5700 33040
rect 122 28041 142 32999
rect 378 28041 5700 32999
rect 5859 32440 5860 33060
rect 6460 32440 6461 33060
rect 5859 32439 6461 32440
rect 5839 31400 6441 31401
rect 5839 30800 5840 31400
rect 6440 30800 6441 31400
rect 5839 30799 6441 30800
rect 122 28000 5700 28041
rect 122 27719 5700 27760
rect 122 22761 142 27719
rect 378 22761 5700 27719
rect 122 22720 5700 22761
rect 122 22439 5700 22480
rect 122 17500 142 22439
rect 100 17481 142 17500
rect 378 17481 5700 22439
rect 100 17440 5700 17481
rect 100 10980 640 17440
rect 100 10660 220 10980
rect 500 10660 640 10980
rect 100 9040 640 10660
rect 100 6840 160 9040
rect 600 6840 640 9040
rect 100 6760 640 6840
rect 6900 6401 7280 33500
rect 19978 19720 22338 19822
rect 19978 17564 20080 19720
rect 22236 17564 22338 19720
rect 19978 8900 22338 17564
rect 19978 6880 20200 8900
rect 22120 6880 22338 8900
rect 19978 6760 22338 6880
rect 6899 6400 7280 6401
rect 6899 6280 6900 6400
rect 7240 6280 7280 6400
rect 6899 6279 7280 6280
rect 6900 5920 7280 6279
rect 6900 5720 7000 5920
rect 7260 5720 7280 5920
rect 6900 5480 7280 5720
rect 6900 5300 6920 5480
rect 7240 5300 7280 5480
rect 6900 5150 7280 5300
rect 17799 5772 23161 5773
rect 17179 3820 17301 3821
rect 17799 3820 17800 5772
rect 17179 3700 17180 3820
rect 17300 3700 17800 3820
rect 17179 3699 17301 3700
rect 6019 3520 6141 3521
rect 6019 3440 6020 3520
rect 6140 3440 6141 3520
rect 6019 3439 6141 3440
rect 6040 3121 6120 3439
rect 5962 3080 12660 3121
rect 5962 2 5982 3080
rect 6218 2 12660 3080
rect 17799 412 17800 3700
rect 23160 412 23161 5772
rect 17799 411 23161 412
rect 17300 140 18080 160
rect 17300 40 17320 140
rect 17420 124 23228 140
rect 17420 60 17748 124
rect 23212 60 23228 124
rect 17420 44 23228 60
rect 17420 40 18080 44
rect 17319 39 17421 40
rect 5962 -39 12660 2
<< via4 >>
rect 142 28041 378 32999
rect 5860 32440 6460 33060
rect 5840 30800 6440 31400
rect 142 22761 378 27719
rect 142 17481 378 22439
rect 20080 17564 22236 19720
rect 11920 3740 12280 3760
rect 11920 3540 11960 3740
rect 11960 3540 12260 3740
rect 12260 3540 12280 3740
rect 11920 3480 12280 3540
rect 5982 2 6218 3080
<< mimcap2 >>
rect 740 32920 5620 32960
rect 740 28120 780 32920
rect 5580 28120 5620 32920
rect 740 28080 5620 28120
rect 740 27640 5620 27680
rect 740 22840 780 27640
rect 5580 22840 5620 27640
rect 740 22800 5620 22840
rect 740 22360 5620 22400
rect 740 17560 780 22360
rect 5580 17560 5620 22360
rect 740 17520 5620 17560
rect 6580 3001 12580 3041
rect 6580 81 6620 3001
rect 12540 81 12580 3001
rect 6580 41 12580 81
<< mimcap2contact >>
rect 780 28120 5580 32920
rect 780 22840 5580 27640
rect 780 17560 5580 22360
rect 6620 81 12540 3001
<< metal5 >>
rect 100 32999 420 33160
rect 100 28041 142 32999
rect 378 28041 420 32999
rect 3020 32944 3340 33160
rect 4939 33060 30680 33122
rect 4939 32944 5860 33060
rect 756 32920 5860 32944
rect 756 28120 780 32920
rect 5580 32440 5860 32920
rect 6460 32440 30680 33060
rect 5580 31400 30680 32440
rect 5580 30800 5840 31400
rect 6440 30800 30680 31400
rect 5580 30760 30680 30800
rect 5580 28120 5604 30760
rect 756 28096 5604 28120
rect 100 27719 420 28041
rect 100 22761 142 27719
rect 378 22761 420 27719
rect 3020 27664 3340 28096
rect 6680 27980 27898 30340
rect 756 27640 5604 27664
rect 756 22840 780 27640
rect 5580 22840 5604 27640
rect 756 22816 5604 22840
rect 100 22439 420 22761
rect 100 17481 142 22439
rect 378 17481 420 22439
rect 3020 22384 3340 22816
rect 756 22360 5604 22384
rect 756 17560 780 22360
rect 5580 17560 5604 22360
rect 756 17536 5604 17560
rect 100 17320 420 17481
rect 3020 17320 3340 17536
rect 6680 11482 9040 27980
rect 9460 25200 25118 27560
rect 9460 14262 11820 25200
rect 12240 22420 22338 24780
rect 12240 17042 14600 22420
rect 19978 19720 22338 22420
rect 19978 17564 20080 19720
rect 22236 17564 22338 19720
rect 19978 17462 22338 17564
rect 22758 17042 25118 25200
rect 12240 14682 25118 17042
rect 25538 14262 27898 27980
rect 9460 11902 27898 14262
rect 28318 11482 30680 30760
rect 6680 9122 30680 11482
rect 11896 3760 12304 3784
rect 11896 3480 11920 3760
rect 12280 3480 12304 3760
rect 11896 3456 12304 3480
rect 5940 3080 6260 3122
rect 5940 2 5982 3080
rect 6218 2 6260 3080
rect 11940 3025 12280 3456
rect 6596 3001 12564 3025
rect 6596 81 6620 3001
rect 12540 81 12564 3001
rect 6596 57 12564 81
rect 5940 -40 6260 2
<< comment >>
rect 6660 6760 6680 6780
<< labels >>
flabel metal1 6040 33620 6240 33820 0 FreeSans 6400 0 0 0 vd
port 0 nsew
flabel metal1 -60 -1180 140 -980 0 FreeSans 6400 0 0 0 gnd
port 1 nsew
flabel metal1 -320 10720 -120 10920 0 FreeSans 6400 0 0 0 out
port 3 nsew
flabel metal1 4680 -1800 4880 -1600 0 FreeSans 6400 0 0 0 ib
port 5 nsew
flabel metal1 14280 -1800 14480 -1600 0 FreeSans 6400 0 0 0 vpwr
port 4 nsew
flabel metal1 13080 -1800 13280 -1600 0 FreeSans 6400 0 0 0 clk
port 2 nsew
flabel metal1 5262 5516 5292 5520 0 FreeSans 1600 0 0 0 vts
flabel metal1 4306 3508 4334 3538 0 FreeSans 1600 0 0 0 vtd
flabel metal1 13376 5282 13494 5370 0 FreeSans 1600 0 0 0 out_buff
flabel metal1 11842 6654 11886 6698 0 FreeSans 800 0 0 0 out_sigma
flabel metal1 6040 33140 6240 33340 0 FreeSans 256 0 0 0 ask-modulator_0.vd
flabel metal1 1040 6560 1240 6760 0 FreeSans 256 0 0 0 ask-modulator_0.gnd
flabel metal1 -80 10720 120 10920 0 FreeSans 256 0 0 0 ask-modulator_0.out
flabel metal1 -80 11260 120 11460 0 FreeSans 256 0 0 0 ask-modulator_0.in
flabel metal1 14300 4140 14500 4340 0 FreeSans 256 0 0 0 sigma-delta_0.in
flabel metal1 14300 2580 14500 2780 0 FreeSans 256 0 0 0 sigma-delta_0.clk
flabel metal1 14300 2020 14500 2220 0 FreeSans 256 0 0 0 sigma-delta_0.reset_b_dff
flabel metal1 15720 0 15920 200 0 FreeSans 256 0 0 0 sigma-delta_0.gnd
flabel metal1 14300 3240 14500 3440 0 FreeSans 256 0 0 0 sigma-delta_0.out
flabel metal1 17340 5680 17540 5880 0 FreeSans 256 0 0 0 sigma-delta_0.vd
flabel metal1 14300 2920 14500 3120 0 FreeSans 256 0 0 0 sigma-delta_0.vpwr
flabel locali 16352 2686 16381 2721 0 FreeSans 200 0 0 0 sigma-delta_0.x1.Q
flabel locali 16654 2689 16676 2722 0 FreeSans 200 0 0 0 sigma-delta_0.x1.Q_N
flabel locali 16079 2621 16113 2655 0 FreeSans 400 0 0 0 sigma-delta_0.x1.RESET_B
flabel locali 14903 2757 14937 2791 0 FreeSans 400 0 0 0 sigma-delta_0.x1.D
flabel locali 14628 2757 14662 2791 0 FreeSans 400 0 0 0 sigma-delta_0.x1.CLK
flabel locali 14628 2689 14662 2723 0 FreeSans 400 0 0 0 sigma-delta_0.x1.CLK
flabel locali 16079 2689 16113 2723 0 FreeSans 400 0 0 0 sigma-delta_0.x1.RESET_B
flabel metal1 14627 2451 14661 2485 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VGND
flabel metal1 14627 2995 14661 3029 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VPWR
flabel nwell 14627 2995 14661 3029 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VPB
flabel pwell 14627 2451 14661 2485 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VNB
rlabel comment 14598 2468 14598 2468 4 sigma-delta_0.x1.dfrbp_1
rlabel locali 16079 2595 16127 2675 1 sigma-delta_0.x1.RESET_B
rlabel locali 16019 2675 16127 2749 1 sigma-delta_0.x1.RESET_B
rlabel metal1 16067 2615 16125 2624 1 sigma-delta_0.x1.RESET_B
rlabel metal1 16007 2661 16065 2724 1 sigma-delta_0.x1.RESET_B
rlabel metal1 16007 2652 16125 2661 1 sigma-delta_0.x1.RESET_B
rlabel metal1 15347 2652 15477 2661 1 sigma-delta_0.x1.RESET_B
rlabel metal1 15347 2624 16125 2652 1 sigma-delta_0.x1.RESET_B
rlabel metal1 15347 2615 15477 2624 1 sigma-delta_0.x1.RESET_B
rlabel metal1 14598 2420 16714 2516 1 sigma-delta_0.x1.VGND
rlabel metal1 14598 2964 16714 3060 1 sigma-delta_0.x1.VPWR
flabel metal1 480 5300 680 5500 0 FreeSans 256 0 0 0 sensor_0.vd
flabel metal1 160 0 360 200 0 FreeSans 256 0 0 0 sensor_0.gnd
flabel metal1 4040 2900 4240 3100 0 FreeSans 256 0 0 0 sensor_0.vts
flabel metal1 4040 3360 4240 3560 0 FreeSans 256 0 0 0 sensor_0.vtd
flabel metal2 860 3580 880 3600 0 FreeSans 800 0 0 0 sensor_0.a
flabel metal2 2380 4440 2400 4460 0 FreeSans 800 0 0 0 sensor_0.d
flabel metal1 2500 3940 2520 3980 0 FreeSans 800 0 0 0 sensor_0.c
flabel metal2 2960 2220 2960 2240 0 FreeSans 800 0 0 0 sensor_0.b
flabel metal1 6280 6240 6480 6440 0 FreeSans 256 0 0 0 buffer_0.vd
flabel metal2 7240 4620 7260 4640 0 FreeSans 800 0 0 0 buffer_0.d
flabel metal1 12600 5220 12800 5420 0 FreeSans 256 0 0 0 buffer_0.out
flabel metal1 5640 5340 5840 5540 0 FreeSans 256 0 0 0 buffer_0.in
flabel metal2 7700 5480 7720 5480 0 FreeSans 800 0 0 0 buffer_0.a
flabel metal2 6720 4620 6740 4640 0 FreeSans 800 0 0 0 buffer_0.c
flabel metal2 10740 5460 10740 5460 0 FreeSans 800 0 0 0 buffer_0.b
flabel metal1 5640 4460 5840 4660 0 FreeSans 256 0 0 0 buffer_0.ib
flabel metal1 5640 3700 5840 3900 0 FreeSans 256 0 0 0 buffer_0.gnd
<< end >>
