magic
tech sky130A
timestamp 1655563127
<< pwell >>
rect -1498 -155 1498 155
<< nmos >>
rect -1400 -50 1400 50
<< ndiff >>
rect -1429 44 -1400 50
rect -1429 -44 -1423 44
rect -1406 -44 -1400 44
rect -1429 -50 -1400 -44
rect 1400 44 1429 50
rect 1400 -44 1406 44
rect 1423 -44 1429 44
rect 1400 -50 1429 -44
<< ndiffc >>
rect -1423 -44 -1406 44
rect 1406 -44 1423 44
<< psubdiff >>
rect -1480 120 -1432 137
rect 1432 120 1480 137
rect -1480 89 -1463 120
rect 1463 89 1480 120
rect -1480 -120 -1463 -89
rect 1463 -120 1480 -89
rect -1480 -137 -1432 -120
rect 1432 -137 1480 -120
<< psubdiffcont >>
rect -1432 120 1432 137
rect -1480 -89 -1463 89
rect 1463 -89 1480 89
rect -1432 -137 1432 -120
<< poly >>
rect -1400 86 1400 94
rect -1400 69 -1392 86
rect 1392 69 1400 86
rect -1400 50 1400 69
rect -1400 -69 1400 -50
rect -1400 -86 -1392 -69
rect 1392 -86 1400 -69
rect -1400 -94 1400 -86
<< polycont >>
rect -1392 69 1392 86
rect -1392 -86 1392 -69
<< locali >>
rect -1480 120 -1432 137
rect 1432 120 1480 137
rect -1480 89 -1463 120
rect 1463 89 1480 120
rect -1400 69 -1392 86
rect 1392 69 1400 86
rect -1423 44 -1406 52
rect -1423 -52 -1406 -44
rect 1406 44 1423 52
rect 1406 -52 1423 -44
rect -1400 -86 -1392 -69
rect 1392 -86 1400 -69
rect -1480 -120 -1463 -89
rect 1463 -120 1480 -89
rect -1480 -137 -1432 -120
rect 1432 -137 1480 -120
<< viali >>
rect -1392 69 1392 86
rect -1423 -44 -1406 44
rect 1406 -44 1423 44
rect -1392 -86 1392 -69
<< metal1 >>
rect -1398 86 1398 89
rect -1398 69 -1392 86
rect 1392 69 1398 86
rect -1398 66 1398 69
rect -1426 44 -1403 50
rect -1426 -44 -1423 44
rect -1406 -44 -1403 44
rect -1426 -50 -1403 -44
rect 1403 44 1426 50
rect 1403 -44 1406 44
rect 1423 -44 1426 44
rect 1403 -50 1426 -44
rect -1398 -69 1398 -66
rect -1398 -86 -1392 -69
rect 1392 -86 1398 -69
rect -1398 -89 1398 -86
<< properties >>
string FIXED_BBOX -1471 -128 1471 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 28.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
