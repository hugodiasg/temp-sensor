magic
tech sky130A
magscale 1 2
timestamp 1661128600
<< nwell >>
rect -1586 -319 1586 319
<< pmos >>
rect -1390 -100 -1190 100
rect -1132 -100 -932 100
rect -874 -100 -674 100
rect -616 -100 -416 100
rect -358 -100 -158 100
rect -100 -100 100 100
rect 158 -100 358 100
rect 416 -100 616 100
rect 674 -100 874 100
rect 932 -100 1132 100
rect 1190 -100 1390 100
<< pdiff >>
rect -1448 88 -1390 100
rect -1448 -88 -1436 88
rect -1402 -88 -1390 88
rect -1448 -100 -1390 -88
rect -1190 88 -1132 100
rect -1190 -88 -1178 88
rect -1144 -88 -1132 88
rect -1190 -100 -1132 -88
rect -932 88 -874 100
rect -932 -88 -920 88
rect -886 -88 -874 88
rect -932 -100 -874 -88
rect -674 88 -616 100
rect -674 -88 -662 88
rect -628 -88 -616 88
rect -674 -100 -616 -88
rect -416 88 -358 100
rect -416 -88 -404 88
rect -370 -88 -358 88
rect -416 -100 -358 -88
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
rect 358 88 416 100
rect 358 -88 370 88
rect 404 -88 416 88
rect 358 -100 416 -88
rect 616 88 674 100
rect 616 -88 628 88
rect 662 -88 674 88
rect 616 -100 674 -88
rect 874 88 932 100
rect 874 -88 886 88
rect 920 -88 932 88
rect 874 -100 932 -88
rect 1132 88 1190 100
rect 1132 -88 1144 88
rect 1178 -88 1190 88
rect 1132 -100 1190 -88
rect 1390 88 1448 100
rect 1390 -88 1402 88
rect 1436 -88 1448 88
rect 1390 -100 1448 -88
<< pdiffc >>
rect -1436 -88 -1402 88
rect -1178 -88 -1144 88
rect -920 -88 -886 88
rect -662 -88 -628 88
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
rect 628 -88 662 88
rect 886 -88 920 88
rect 1144 -88 1178 88
rect 1402 -88 1436 88
<< nsubdiff >>
rect -1550 249 -1454 283
rect 1454 249 1550 283
rect -1550 187 -1516 249
rect 1516 187 1550 249
rect -1550 -249 -1516 -187
rect 1516 -249 1550 -187
rect -1550 -283 -1454 -249
rect 1454 -283 1550 -249
<< nsubdiffcont >>
rect -1454 249 1454 283
rect -1550 -187 -1516 187
rect 1516 -187 1550 187
rect -1454 -283 1454 -249
<< poly >>
rect -1390 181 -1190 197
rect -1390 147 -1374 181
rect -1206 147 -1190 181
rect -1390 100 -1190 147
rect -1132 181 -932 197
rect -1132 147 -1116 181
rect -948 147 -932 181
rect -1132 100 -932 147
rect -874 181 -674 197
rect -874 147 -858 181
rect -690 147 -674 181
rect -874 100 -674 147
rect -616 181 -416 197
rect -616 147 -600 181
rect -432 147 -416 181
rect -616 100 -416 147
rect -358 181 -158 197
rect -358 147 -342 181
rect -174 147 -158 181
rect -358 100 -158 147
rect -100 181 100 197
rect -100 147 -84 181
rect 84 147 100 181
rect -100 100 100 147
rect 158 181 358 197
rect 158 147 174 181
rect 342 147 358 181
rect 158 100 358 147
rect 416 181 616 197
rect 416 147 432 181
rect 600 147 616 181
rect 416 100 616 147
rect 674 181 874 197
rect 674 147 690 181
rect 858 147 874 181
rect 674 100 874 147
rect 932 181 1132 197
rect 932 147 948 181
rect 1116 147 1132 181
rect 932 100 1132 147
rect 1190 181 1390 197
rect 1190 147 1206 181
rect 1374 147 1390 181
rect 1190 100 1390 147
rect -1390 -147 -1190 -100
rect -1390 -181 -1374 -147
rect -1206 -181 -1190 -147
rect -1390 -197 -1190 -181
rect -1132 -147 -932 -100
rect -1132 -181 -1116 -147
rect -948 -181 -932 -147
rect -1132 -197 -932 -181
rect -874 -147 -674 -100
rect -874 -181 -858 -147
rect -690 -181 -674 -147
rect -874 -197 -674 -181
rect -616 -147 -416 -100
rect -616 -181 -600 -147
rect -432 -181 -416 -147
rect -616 -197 -416 -181
rect -358 -147 -158 -100
rect -358 -181 -342 -147
rect -174 -181 -158 -147
rect -358 -197 -158 -181
rect -100 -147 100 -100
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -100 -197 100 -181
rect 158 -147 358 -100
rect 158 -181 174 -147
rect 342 -181 358 -147
rect 158 -197 358 -181
rect 416 -147 616 -100
rect 416 -181 432 -147
rect 600 -181 616 -147
rect 416 -197 616 -181
rect 674 -147 874 -100
rect 674 -181 690 -147
rect 858 -181 874 -147
rect 674 -197 874 -181
rect 932 -147 1132 -100
rect 932 -181 948 -147
rect 1116 -181 1132 -147
rect 932 -197 1132 -181
rect 1190 -147 1390 -100
rect 1190 -181 1206 -147
rect 1374 -181 1390 -147
rect 1190 -197 1390 -181
<< polycont >>
rect -1374 147 -1206 181
rect -1116 147 -948 181
rect -858 147 -690 181
rect -600 147 -432 181
rect -342 147 -174 181
rect -84 147 84 181
rect 174 147 342 181
rect 432 147 600 181
rect 690 147 858 181
rect 948 147 1116 181
rect 1206 147 1374 181
rect -1374 -181 -1206 -147
rect -1116 -181 -948 -147
rect -858 -181 -690 -147
rect -600 -181 -432 -147
rect -342 -181 -174 -147
rect -84 -181 84 -147
rect 174 -181 342 -147
rect 432 -181 600 -147
rect 690 -181 858 -147
rect 948 -181 1116 -147
rect 1206 -181 1374 -147
<< locali >>
rect -1550 249 -1454 283
rect 1454 249 1550 283
rect -1550 187 -1516 249
rect 1516 187 1550 249
rect -1390 147 -1374 181
rect -1206 147 -1190 181
rect -1132 147 -1116 181
rect -948 147 -932 181
rect -874 147 -858 181
rect -690 147 -674 181
rect -616 147 -600 181
rect -432 147 -416 181
rect -358 147 -342 181
rect -174 147 -158 181
rect -100 147 -84 181
rect 84 147 100 181
rect 158 147 174 181
rect 342 147 358 181
rect 416 147 432 181
rect 600 147 616 181
rect 674 147 690 181
rect 858 147 874 181
rect 932 147 948 181
rect 1116 147 1132 181
rect 1190 147 1206 181
rect 1374 147 1390 181
rect -1436 88 -1402 104
rect -1436 -104 -1402 -88
rect -1178 88 -1144 104
rect -1178 -104 -1144 -88
rect -920 88 -886 104
rect -920 -104 -886 -88
rect -662 88 -628 104
rect -662 -104 -628 -88
rect -404 88 -370 104
rect -404 -104 -370 -88
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect 370 88 404 104
rect 370 -104 404 -88
rect 628 88 662 104
rect 628 -104 662 -88
rect 886 88 920 104
rect 886 -104 920 -88
rect 1144 88 1178 104
rect 1144 -104 1178 -88
rect 1402 88 1436 104
rect 1402 -104 1436 -88
rect -1390 -181 -1374 -147
rect -1206 -181 -1190 -147
rect -1132 -181 -1116 -147
rect -948 -181 -932 -147
rect -874 -181 -858 -147
rect -690 -181 -674 -147
rect -616 -181 -600 -147
rect -432 -181 -416 -147
rect -358 -181 -342 -147
rect -174 -181 -158 -147
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect 158 -181 174 -147
rect 342 -181 358 -147
rect 416 -181 432 -147
rect 600 -181 616 -147
rect 674 -181 690 -147
rect 858 -181 874 -147
rect 932 -181 948 -147
rect 1116 -181 1132 -147
rect 1190 -181 1206 -147
rect 1374 -181 1390 -147
rect -1550 -249 -1516 -187
rect 1516 -249 1550 -187
rect -1550 -283 -1454 -249
rect 1454 -283 1550 -249
<< viali >>
rect -1374 147 -1206 181
rect -1116 147 -948 181
rect -858 147 -690 181
rect -600 147 -432 181
rect -342 147 -174 181
rect -84 147 84 181
rect 174 147 342 181
rect 432 147 600 181
rect 690 147 858 181
rect 948 147 1116 181
rect 1206 147 1374 181
rect -1436 -88 -1402 88
rect -1178 -88 -1144 88
rect -920 -88 -886 88
rect -662 -88 -628 88
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
rect 628 -88 662 88
rect 886 -88 920 88
rect 1144 -88 1178 88
rect 1402 -88 1436 88
rect -1374 -181 -1206 -147
rect -1116 -181 -948 -147
rect -858 -181 -690 -147
rect -600 -181 -432 -147
rect -342 -181 -174 -147
rect -84 -181 84 -147
rect 174 -181 342 -147
rect 432 -181 600 -147
rect 690 -181 858 -147
rect 948 -181 1116 -147
rect 1206 -181 1374 -147
<< metal1 >>
rect -1386 181 -1194 187
rect -1386 147 -1374 181
rect -1206 147 -1194 181
rect -1386 141 -1194 147
rect -1128 181 -936 187
rect -1128 147 -1116 181
rect -948 147 -936 181
rect -1128 141 -936 147
rect -870 181 -678 187
rect -870 147 -858 181
rect -690 147 -678 181
rect -870 141 -678 147
rect -612 181 -420 187
rect -612 147 -600 181
rect -432 147 -420 181
rect -612 141 -420 147
rect -354 181 -162 187
rect -354 147 -342 181
rect -174 147 -162 181
rect -354 141 -162 147
rect -96 181 96 187
rect -96 147 -84 181
rect 84 147 96 181
rect -96 141 96 147
rect 162 181 354 187
rect 162 147 174 181
rect 342 147 354 181
rect 162 141 354 147
rect 420 181 612 187
rect 420 147 432 181
rect 600 147 612 181
rect 420 141 612 147
rect 678 181 870 187
rect 678 147 690 181
rect 858 147 870 181
rect 678 141 870 147
rect 936 181 1128 187
rect 936 147 948 181
rect 1116 147 1128 181
rect 936 141 1128 147
rect 1194 181 1386 187
rect 1194 147 1206 181
rect 1374 147 1386 181
rect 1194 141 1386 147
rect -1442 88 -1396 100
rect -1442 -88 -1436 88
rect -1402 -88 -1396 88
rect -1442 -100 -1396 -88
rect -1184 88 -1138 100
rect -1184 -88 -1178 88
rect -1144 -88 -1138 88
rect -1184 -100 -1138 -88
rect -926 88 -880 100
rect -926 -88 -920 88
rect -886 -88 -880 88
rect -926 -100 -880 -88
rect -668 88 -622 100
rect -668 -88 -662 88
rect -628 -88 -622 88
rect -668 -100 -622 -88
rect -410 88 -364 100
rect -410 -88 -404 88
rect -370 -88 -364 88
rect -410 -100 -364 -88
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect 364 88 410 100
rect 364 -88 370 88
rect 404 -88 410 88
rect 364 -100 410 -88
rect 622 88 668 100
rect 622 -88 628 88
rect 662 -88 668 88
rect 622 -100 668 -88
rect 880 88 926 100
rect 880 -88 886 88
rect 920 -88 926 88
rect 880 -100 926 -88
rect 1138 88 1184 100
rect 1138 -88 1144 88
rect 1178 -88 1184 88
rect 1138 -100 1184 -88
rect 1396 88 1442 100
rect 1396 -88 1402 88
rect 1436 -88 1442 88
rect 1396 -100 1442 -88
rect -1386 -147 -1194 -141
rect -1386 -181 -1374 -147
rect -1206 -181 -1194 -147
rect -1386 -187 -1194 -181
rect -1128 -147 -936 -141
rect -1128 -181 -1116 -147
rect -948 -181 -936 -147
rect -1128 -187 -936 -181
rect -870 -147 -678 -141
rect -870 -181 -858 -147
rect -690 -181 -678 -147
rect -870 -187 -678 -181
rect -612 -147 -420 -141
rect -612 -181 -600 -147
rect -432 -181 -420 -147
rect -612 -187 -420 -181
rect -354 -147 -162 -141
rect -354 -181 -342 -147
rect -174 -181 -162 -147
rect -354 -187 -162 -181
rect -96 -147 96 -141
rect -96 -181 -84 -147
rect 84 -181 96 -147
rect -96 -187 96 -181
rect 162 -147 354 -141
rect 162 -181 174 -147
rect 342 -181 354 -147
rect 162 -187 354 -181
rect 420 -147 612 -141
rect 420 -181 432 -147
rect 600 -181 612 -147
rect 420 -187 612 -181
rect 678 -147 870 -141
rect 678 -181 690 -147
rect 858 -181 870 -147
rect 678 -187 870 -181
rect 936 -147 1128 -141
rect 936 -181 948 -147
rect 1116 -181 1128 -147
rect 936 -187 1128 -181
rect 1194 -147 1386 -141
rect 1194 -181 1206 -147
rect 1374 -181 1386 -147
rect 1194 -187 1386 -181
<< properties >>
string FIXED_BBOX -1533 -266 1533 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
