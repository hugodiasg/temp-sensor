magic
tech sky130A
timestamp 1700075225
<< pwell >>
rect -1798 -155 1798 155
<< nmos >>
rect -1700 -50 1700 50
<< ndiff >>
rect -1729 44 -1700 50
rect -1729 -44 -1723 44
rect -1706 -44 -1700 44
rect -1729 -50 -1700 -44
rect 1700 44 1729 50
rect 1700 -44 1706 44
rect 1723 -44 1729 44
rect 1700 -50 1729 -44
<< ndiffc >>
rect -1723 -44 -1706 44
rect 1706 -44 1723 44
<< psubdiff >>
rect -1780 120 -1732 137
rect 1732 120 1780 137
rect -1780 89 -1763 120
rect 1763 89 1780 120
rect -1780 -120 -1763 -89
rect 1763 -120 1780 -89
rect -1780 -137 -1732 -120
rect 1732 -137 1780 -120
<< psubdiffcont >>
rect -1732 120 1732 137
rect -1780 -89 -1763 89
rect 1763 -89 1780 89
rect -1732 -137 1732 -120
<< poly >>
rect -1700 86 1700 94
rect -1700 69 -1692 86
rect 1692 69 1700 86
rect -1700 50 1700 69
rect -1700 -69 1700 -50
rect -1700 -86 -1692 -69
rect 1692 -86 1700 -69
rect -1700 -94 1700 -86
<< polycont >>
rect -1692 69 1692 86
rect -1692 -86 1692 -69
<< locali >>
rect -1780 120 -1732 137
rect 1732 120 1780 137
rect -1780 89 -1763 120
rect 1763 89 1780 120
rect -1700 69 -1692 86
rect 1692 69 1700 86
rect -1723 44 -1706 52
rect -1723 -52 -1706 -44
rect 1706 44 1723 52
rect 1706 -52 1723 -44
rect -1700 -86 -1692 -69
rect 1692 -86 1700 -69
rect -1780 -120 -1763 -89
rect 1763 -120 1780 -89
rect -1780 -137 -1732 -120
rect 1732 -137 1780 -120
<< viali >>
rect -1692 69 1692 86
rect -1723 -44 -1706 44
rect 1706 -44 1723 44
rect -1692 -86 1692 -69
<< metal1 >>
rect -1698 86 1698 89
rect -1698 69 -1692 86
rect 1692 69 1698 86
rect -1698 66 1698 69
rect -1726 44 -1703 50
rect -1726 -44 -1723 44
rect -1706 -44 -1703 44
rect -1726 -50 -1703 -44
rect 1703 44 1726 50
rect 1703 -44 1706 44
rect 1723 -44 1726 44
rect 1703 -50 1726 -44
rect -1698 -69 1698 -66
rect -1698 -86 -1692 -69
rect 1692 -86 1698 -69
rect -1698 -89 1698 -86
<< properties >>
string FIXED_BBOX -1771 -128 1771 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 34 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
