magic
tech sky130A
timestamp 1700075225
<< pwell >>
rect -1698 -155 1698 155
<< nmos >>
rect -1600 -50 1600 50
<< ndiff >>
rect -1629 44 -1600 50
rect -1629 -44 -1623 44
rect -1606 -44 -1600 44
rect -1629 -50 -1600 -44
rect 1600 44 1629 50
rect 1600 -44 1606 44
rect 1623 -44 1629 44
rect 1600 -50 1629 -44
<< ndiffc >>
rect -1623 -44 -1606 44
rect 1606 -44 1623 44
<< psubdiff >>
rect -1680 120 -1632 137
rect 1632 120 1680 137
rect -1680 89 -1663 120
rect 1663 89 1680 120
rect -1680 -120 -1663 -89
rect 1663 -120 1680 -89
rect -1680 -137 -1632 -120
rect 1632 -137 1680 -120
<< psubdiffcont >>
rect -1632 120 1632 137
rect -1680 -89 -1663 89
rect 1663 -89 1680 89
rect -1632 -137 1632 -120
<< poly >>
rect -1600 86 1600 94
rect -1600 69 -1592 86
rect 1592 69 1600 86
rect -1600 50 1600 69
rect -1600 -69 1600 -50
rect -1600 -86 -1592 -69
rect 1592 -86 1600 -69
rect -1600 -94 1600 -86
<< polycont >>
rect -1592 69 1592 86
rect -1592 -86 1592 -69
<< locali >>
rect -1680 120 -1632 137
rect 1632 120 1680 137
rect -1680 89 -1663 120
rect 1663 89 1680 120
rect -1600 69 -1592 86
rect 1592 69 1600 86
rect -1623 44 -1606 52
rect -1623 -52 -1606 -44
rect 1606 44 1623 52
rect 1606 -52 1623 -44
rect -1600 -86 -1592 -69
rect 1592 -86 1600 -69
rect -1680 -120 -1663 -89
rect 1663 -120 1680 -89
rect -1680 -137 -1632 -120
rect 1632 -137 1680 -120
<< viali >>
rect -1592 69 1592 86
rect -1623 -44 -1606 44
rect 1606 -44 1623 44
rect -1592 -86 1592 -69
<< metal1 >>
rect -1598 86 1598 89
rect -1598 69 -1592 86
rect 1592 69 1598 86
rect -1598 66 1598 69
rect -1626 44 -1603 50
rect -1626 -44 -1623 44
rect -1606 -44 -1603 44
rect -1626 -50 -1603 -44
rect 1603 44 1626 50
rect 1603 -44 1606 44
rect 1623 -44 1626 44
rect 1603 -50 1626 -44
rect -1598 -69 1598 -66
rect -1598 -86 -1592 -69
rect 1592 -86 1598 -69
rect -1598 -89 1598 -86
<< properties >>
string FIXED_BBOX -1671 -128 1671 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 32 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
