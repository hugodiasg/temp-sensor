** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/nmos_tb.sch
**.subckt nmos_tb
Va in GND 1.8
V2 out GND 3.3
XM1 out in GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=21 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.dc V2 0V 5 0.01V
.control
run
plot -I(v2)
plot out/(-i(v2))
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
