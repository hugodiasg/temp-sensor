magic
tech sky130A
magscale 1 2
timestamp 1645799446
<< metal4 >>
rect -2622 10281 2622 10322
rect -2622 5277 2366 10281
rect 2602 5277 2622 10281
rect -2622 5236 2622 5277
rect -2622 5095 2622 5136
rect -2622 91 2366 5095
rect 2602 91 2622 5095
rect -2622 50 2622 91
rect -2622 -91 2622 -50
rect -2622 -5095 2366 -91
rect 2602 -5095 2622 -91
rect -2622 -5136 2622 -5095
rect -2622 -5277 2622 -5236
rect -2622 -10281 2366 -5277
rect 2602 -10281 2622 -5277
rect -2622 -10322 2622 -10281
<< via4 >>
rect 2366 5277 2602 10281
rect 2366 91 2602 5095
rect 2366 -5095 2602 -91
rect 2366 -10281 2602 -5277
<< mimcap2 >>
rect -2522 10182 2364 10222
rect -2522 5376 -2001 10182
rect 1843 5376 2364 10182
rect -2522 5336 2364 5376
rect -2522 4996 2364 5036
rect -2522 190 -2001 4996
rect 1843 190 2364 4996
rect -2522 150 2364 190
rect -2522 -190 2364 -150
rect -2522 -4996 -2001 -190
rect 1843 -4996 2364 -190
rect -2522 -5036 2364 -4996
rect -2522 -5376 2364 -5336
rect -2522 -10182 -2001 -5376
rect 1843 -10182 2364 -5376
rect -2522 -10222 2364 -10182
<< mimcap2contact >>
rect -2001 5376 1843 10182
rect -2001 190 1843 4996
rect -2001 -4996 1843 -190
rect -2001 -10182 1843 -5376
<< metal5 >>
rect -239 10206 81 10372
rect 2324 10281 2644 10372
rect -2025 10182 1867 10206
rect -2025 5376 -2001 10182
rect 1843 5376 1867 10182
rect -2025 5352 1867 5376
rect -239 5020 81 5352
rect 2324 5277 2366 10281
rect 2602 5277 2644 10281
rect 2324 5095 2644 5277
rect -2025 4996 1867 5020
rect -2025 190 -2001 4996
rect 1843 190 1867 4996
rect -2025 166 1867 190
rect -239 -166 81 166
rect 2324 91 2366 5095
rect 2602 91 2644 5095
rect 2324 -91 2644 91
rect -2025 -190 1867 -166
rect -2025 -4996 -2001 -190
rect 1843 -4996 1867 -190
rect -2025 -5020 1867 -4996
rect -239 -5352 81 -5020
rect 2324 -5095 2366 -91
rect 2602 -5095 2644 -91
rect 2324 -5277 2644 -5095
rect -2025 -5376 1867 -5352
rect -2025 -10182 -2001 -5376
rect 1843 -10182 1867 -5376
rect -2025 -10206 1867 -10182
rect -239 -10372 81 -10206
rect 2324 -10281 2366 -5277
rect 2602 -10281 2644 -5277
rect 2324 -10372 2644 -10281
<< properties >>
string FIXED_BBOX -2622 5236 2464 10322
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.43 l 24.43 val 1.212k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
