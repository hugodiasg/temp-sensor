magic
tech sky130A
magscale 1 2
timestamp 1644351742
<< metal4 >>
rect -2459 7199 2459 7240
rect -2459 2521 2203 7199
rect 2439 2521 2459 7199
rect -2459 2480 2459 2521
rect -2459 2339 2459 2380
rect -2459 -2339 2203 2339
rect 2439 -2339 2459 2339
rect -2459 -2380 2459 -2339
rect -2459 -2521 2459 -2480
rect -2459 -7199 2203 -2521
rect 2439 -7199 2459 -2521
rect -2459 -7240 2459 -7199
<< via4 >>
rect 2203 2521 2439 7199
rect 2203 -2339 2439 2339
rect 2203 -7199 2439 -2521
<< mimcap2 >>
rect -2359 7100 2201 7140
rect -2359 2620 -1871 7100
rect 1713 2620 2201 7100
rect -2359 2580 2201 2620
rect -2359 2240 2201 2280
rect -2359 -2240 -1871 2240
rect 1713 -2240 2201 2240
rect -2359 -2280 2201 -2240
rect -2359 -2620 2201 -2580
rect -2359 -7100 -1871 -2620
rect 1713 -7100 2201 -2620
rect -2359 -7140 2201 -7100
<< mimcap2contact >>
rect -1871 2620 1713 7100
rect -1871 -2240 1713 2240
rect -1871 -7100 1713 -2620
<< metal5 >>
rect -239 7124 81 7290
rect 2161 7199 2481 7290
rect -1895 7100 1737 7124
rect -1895 2620 -1871 7100
rect 1713 2620 1737 7100
rect -1895 2596 1737 2620
rect -239 2264 81 2596
rect 2161 2521 2203 7199
rect 2439 2521 2481 7199
rect 2161 2339 2481 2521
rect -1895 2240 1737 2264
rect -1895 -2240 -1871 2240
rect 1713 -2240 1737 2240
rect -1895 -2264 1737 -2240
rect -239 -2596 81 -2264
rect 2161 -2339 2203 2339
rect 2439 -2339 2481 2339
rect 2161 -2521 2481 -2339
rect -1895 -2620 1737 -2596
rect -1895 -7100 -1871 -2620
rect 1713 -7100 1737 -2620
rect -1895 -7124 1737 -7100
rect -239 -7290 81 -7124
rect 2161 -7199 2203 -2521
rect 2439 -7199 2481 -2521
rect 2161 -7290 2481 -7199
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2459 2480 2301 7240
string parameters w 22.8 l 22.8 val 1.057k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
