magic
tech sky130A
magscale 1 2
timestamp 1645495691
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
use sky130_fd_pr__cap_mim_m3_2_L3GQVG  XC0
timestamp 1645495691
transform 1 0 6819 0 1 50633
box -2635 -7818 2657 7818
use sky130_fd_pr__cap_mim_m3_2_H8XJTH  XC1
timestamp 1645495691
transform 1 0 25880 0 1 74404
box -3080 -12204 3102 12204
use l0  l0_0
timestamp 1645495691
transform 1 0 -10799 0 1 -10000
box 32199 32200 70200 71480
use sky130_fd_pr__cap_mim_m3_2_H8XJTH  sky130_fd_pr__cap_mim_m3_2_H8XJTH_0
timestamp 1645495691
transform 1 0 32280 0 1 74404
box -3080 -12204 3102 12204
use sky130_fd_pr__cap_mim_m3_2_H8XJTH  sky130_fd_pr__cap_mim_m3_2_H8XJTH_1
timestamp 1645495691
transform 1 0 38680 0 1 74404
box -3080 -12204 3102 12204
use sky130_fd_pr__cap_mim_m3_2_H8XJTH  sky130_fd_pr__cap_mim_m3_2_H8XJTH_2
timestamp 1645495691
transform 1 0 45080 0 1 74404
box -3080 -12204 3102 12204
use sky130_fd_pr__cap_mim_m3_2_L3GQVG  sky130_fd_pr__cap_mim_m3_2_L3GQVG_0
timestamp 1645495691
transform 1 0 12435 0 1 50618
box -2635 -7818 2657 7818
use sky130_fd_pr__cap_mim_m3_2_L3GQVG  sky130_fd_pr__cap_mim_m3_2_L3GQVG_1
timestamp 1645495691
transform 1 0 18035 0 1 50618
box -2635 -7818 2657 7818
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 128 0 0 0 gnd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 128 0 0 0 out
port 2 nsew
<< end >>
