magic
tech sky130A
magscale 1 2
timestamp 1644351742
<< error_p >>
rect 1837 2596 1845 7124
rect 2157 2521 2165 7199
rect 2477 2479 2485 2701
rect 1837 -2264 1845 2264
rect 2157 -2339 2165 2339
rect 2477 2159 2485 2381
rect 2477 -2381 2485 -2159
rect 1837 -7124 1845 -2596
rect 2157 -7199 2165 -2521
rect 2477 -2701 2485 -2479
<< metal4 >>
rect -2463 7199 2463 7240
rect -2463 2521 2207 7199
rect 2443 2521 2463 7199
rect -2463 2480 2463 2521
rect -2463 2339 2463 2380
rect -2463 -2339 2207 2339
rect 2443 -2339 2463 2339
rect -2463 -2380 2463 -2339
rect -2463 -2521 2463 -2480
rect -2463 -7199 2207 -2521
rect 2443 -7199 2463 -2521
rect -2463 -7240 2463 -7199
<< via4 >>
rect 2207 2521 2443 7199
rect 2207 -2339 2443 2339
rect 2207 -7199 2443 -2521
<< mimcap2 >>
rect -2363 7100 2197 7140
rect -2363 2620 -1987 7100
rect 1821 2620 2197 7100
rect -2363 2580 2197 2620
rect -2363 2240 2197 2280
rect -2363 -2240 -1987 2240
rect 1821 -2240 2197 2240
rect -2363 -2280 2197 -2240
rect -2363 -2620 2197 -2580
rect -2363 -7100 -1987 -2620
rect 1821 -7100 2197 -2620
rect -2363 -7140 2197 -7100
<< mimcap2contact >>
rect -1987 2620 1821 7100
rect -1987 -2240 1821 2240
rect -1987 -7100 1821 -2620
<< metal5 >>
rect -243 7124 77 7290
rect 2157 7241 2477 7290
rect 2157 7199 2485 7241
rect -2011 7100 1845 7124
rect -2011 2620 -1987 7100
rect 1821 2620 1845 7100
rect -2011 2596 1845 2620
rect -243 2264 77 2596
rect 2157 2521 2207 7199
rect 2443 2521 2485 7199
rect 2157 2479 2485 2521
rect 2157 2381 2477 2479
rect 2157 2339 2485 2381
rect -2011 2240 1845 2264
rect -2011 -2240 -1987 2240
rect 1821 -2240 1845 2240
rect -2011 -2264 1845 -2240
rect -243 -2596 77 -2264
rect 2157 -2339 2207 2339
rect 2443 -2339 2485 2339
rect 2157 -2381 2485 -2339
rect 2157 -2479 2477 -2381
rect 2157 -2521 2485 -2479
rect -2011 -2620 1845 -2596
rect -2011 -7100 -1987 -2620
rect 1821 -7100 1845 -2620
rect -2011 -7124 1845 -7100
rect -243 -7290 77 -7124
rect 2157 -7199 2207 -2521
rect 2443 -7199 2485 -2521
rect 2157 -7241 2485 -7199
rect 2157 -7290 2477 -7241
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2463 2480 2297 7240
string parameters w 22.8 l 22.8 val 1.057k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 85
string library sky130
<< end >>
