magic
tech sky130A
magscale 1 2
timestamp 1707923906
<< metal3 >>
rect -2636 7652 2636 7680
rect -2636 2748 2552 7652
rect 2616 2748 2636 7652
rect -2636 2720 2636 2748
rect -2636 2452 2636 2480
rect -2636 -2452 2552 2452
rect 2616 -2452 2636 2452
rect -2636 -2480 2636 -2452
rect -2636 -2748 2636 -2720
rect -2636 -7652 2552 -2748
rect 2616 -7652 2636 -2748
rect -2636 -7680 2636 -7652
<< via3 >>
rect 2552 2748 2616 7652
rect 2552 -2452 2616 2452
rect 2552 -7652 2616 -2748
<< mimcap >>
rect -2596 7600 2304 7640
rect -2596 2800 -2556 7600
rect 2264 2800 2304 7600
rect -2596 2760 2304 2800
rect -2596 2400 2304 2440
rect -2596 -2400 -2556 2400
rect 2264 -2400 2304 2400
rect -2596 -2440 2304 -2400
rect -2596 -2800 2304 -2760
rect -2596 -7600 -2556 -2800
rect 2264 -7600 2304 -2800
rect -2596 -7640 2304 -7600
<< mimcapcontact >>
rect -2556 2800 2264 7600
rect -2556 -2400 2264 2400
rect -2556 -7600 2264 -2800
<< metal4 >>
rect -198 7601 -94 7800
rect 2532 7652 2636 7800
rect -2557 7600 2265 7601
rect -2557 2800 -2556 7600
rect 2264 2800 2265 7600
rect -2557 2799 2265 2800
rect -198 2401 -94 2799
rect 2532 2748 2552 7652
rect 2616 2748 2636 7652
rect 2532 2452 2636 2748
rect -2557 2400 2265 2401
rect -2557 -2400 -2556 2400
rect 2264 -2400 2265 2400
rect -2557 -2401 2265 -2400
rect -198 -2799 -94 -2401
rect 2532 -2452 2552 2452
rect 2616 -2452 2636 2452
rect 2532 -2748 2636 -2452
rect -2557 -2800 2265 -2799
rect -2557 -7600 -2556 -2800
rect 2264 -7600 2265 -2800
rect -2557 -7601 2265 -7600
rect -198 -7800 -94 -7601
rect 2532 -7652 2552 -2748
rect 2616 -7652 2636 -2748
rect 2532 -7800 2636 -7652
<< properties >>
string FIXED_BBOX -2636 2720 2344 7680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 24.5 l 24.4 val 1.214k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
