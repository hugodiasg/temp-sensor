magic
tech sky130A
magscale 1 2
timestamp 1645556896
<< metal4 >>
rect -1200 2980 3000 3000
rect -1200 1820 1796 2980
rect 2956 1820 3000 2980
rect -1200 1800 3000 1820
rect 1793 1795 2998 1800
<< via4 >>
rect 1796 1820 2956 2980
<< metal5 >>
rect 0 28800 30000 30000
rect 0 27000 28200 28200
rect 0 1200 1200 27000
rect 1785 3004 2998 3007
rect 1772 3000 2998 3004
rect 27000 3000 28200 27000
rect 1772 2980 28200 3000
rect 1772 1820 1796 2980
rect 2956 1820 28200 2980
rect 1772 1800 28200 1820
rect 1772 1796 2998 1800
rect 1785 1792 2998 1796
rect 28800 1200 30000 28800
rect 0 0 30000 1200
<< end >>
