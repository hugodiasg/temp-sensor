magic
tech sky130A
magscale 1 2
timestamp 1675569099
<< metal4 >>
rect -12345 10639 -7727 10680
rect -12345 6641 -7983 10639
rect -7747 6641 -7727 10639
rect -12345 6600 -7727 6641
rect -7327 10639 -2709 10680
rect -7327 6641 -2965 10639
rect -2729 6641 -2709 10639
rect -7327 6600 -2709 6641
rect -2309 10639 2309 10680
rect -2309 6641 2053 10639
rect 2289 6641 2309 10639
rect -2309 6600 2309 6641
rect 2709 10639 7327 10680
rect 2709 6641 7071 10639
rect 7307 6641 7327 10639
rect 2709 6600 7327 6641
rect 7727 10639 12345 10680
rect 7727 6641 12089 10639
rect 12325 6641 12345 10639
rect 7727 6600 12345 6641
rect -12345 6319 -7727 6360
rect -12345 2321 -7983 6319
rect -7747 2321 -7727 6319
rect -12345 2280 -7727 2321
rect -7327 6319 -2709 6360
rect -7327 2321 -2965 6319
rect -2729 2321 -2709 6319
rect -7327 2280 -2709 2321
rect -2309 6319 2309 6360
rect -2309 2321 2053 6319
rect 2289 2321 2309 6319
rect -2309 2280 2309 2321
rect 2709 6319 7327 6360
rect 2709 2321 7071 6319
rect 7307 2321 7327 6319
rect 2709 2280 7327 2321
rect 7727 6319 12345 6360
rect 7727 2321 12089 6319
rect 12325 2321 12345 6319
rect 7727 2280 12345 2321
rect -12345 1999 -7727 2040
rect -12345 -1999 -7983 1999
rect -7747 -1999 -7727 1999
rect -12345 -2040 -7727 -1999
rect -7327 1999 -2709 2040
rect -7327 -1999 -2965 1999
rect -2729 -1999 -2709 1999
rect -7327 -2040 -2709 -1999
rect -2309 1999 2309 2040
rect -2309 -1999 2053 1999
rect 2289 -1999 2309 1999
rect -2309 -2040 2309 -1999
rect 2709 1999 7327 2040
rect 2709 -1999 7071 1999
rect 7307 -1999 7327 1999
rect 2709 -2040 7327 -1999
rect 7727 1999 12345 2040
rect 7727 -1999 12089 1999
rect 12325 -1999 12345 1999
rect 7727 -2040 12345 -1999
rect -12345 -2321 -7727 -2280
rect -12345 -6319 -7983 -2321
rect -7747 -6319 -7727 -2321
rect -12345 -6360 -7727 -6319
rect -7327 -2321 -2709 -2280
rect -7327 -6319 -2965 -2321
rect -2729 -6319 -2709 -2321
rect -7327 -6360 -2709 -6319
rect -2309 -2321 2309 -2280
rect -2309 -6319 2053 -2321
rect 2289 -6319 2309 -2321
rect -2309 -6360 2309 -6319
rect 2709 -2321 7327 -2280
rect 2709 -6319 7071 -2321
rect 7307 -6319 7327 -2321
rect 2709 -6360 7327 -6319
rect 7727 -2321 12345 -2280
rect 7727 -6319 12089 -2321
rect 12325 -6319 12345 -2321
rect 7727 -6360 12345 -6319
rect -12345 -6641 -7727 -6600
rect -12345 -10639 -7983 -6641
rect -7747 -10639 -7727 -6641
rect -12345 -10680 -7727 -10639
rect -7327 -6641 -2709 -6600
rect -7327 -10639 -2965 -6641
rect -2729 -10639 -2709 -6641
rect -7327 -10680 -2709 -10639
rect -2309 -6641 2309 -6600
rect -2309 -10639 2053 -6641
rect 2289 -10639 2309 -6641
rect -2309 -10680 2309 -10639
rect 2709 -6641 7327 -6600
rect 2709 -10639 7071 -6641
rect 7307 -10639 7327 -6641
rect 2709 -10680 7327 -10639
rect 7727 -6641 12345 -6600
rect 7727 -10639 12089 -6641
rect 12325 -10639 12345 -6641
rect 7727 -10680 12345 -10639
<< via4 >>
rect -7983 6641 -7747 10639
rect -2965 6641 -2729 10639
rect 2053 6641 2289 10639
rect 7071 6641 7307 10639
rect 12089 6641 12325 10639
rect -7983 2321 -7747 6319
rect -2965 2321 -2729 6319
rect 2053 2321 2289 6319
rect 7071 2321 7307 6319
rect 12089 2321 12325 6319
rect -7983 -1999 -7747 1999
rect -2965 -1999 -2729 1999
rect 2053 -1999 2289 1999
rect 7071 -1999 7307 1999
rect 12089 -1999 12325 1999
rect -7983 -6319 -7747 -2321
rect -2965 -6319 -2729 -2321
rect 2053 -6319 2289 -2321
rect 7071 -6319 7307 -2321
rect 12089 -6319 12325 -2321
rect -7983 -10639 -7747 -6641
rect -2965 -10639 -2729 -6641
rect 2053 -10639 2289 -6641
rect 7071 -10639 7307 -6641
rect 12089 -10639 12325 -6641
<< mimcap2 >>
rect -12265 10560 -8345 10600
rect -12265 6720 -12225 10560
rect -8385 6720 -8345 10560
rect -12265 6680 -8345 6720
rect -7247 10560 -3327 10600
rect -7247 6720 -7207 10560
rect -3367 6720 -3327 10560
rect -7247 6680 -3327 6720
rect -2229 10560 1691 10600
rect -2229 6720 -2189 10560
rect 1651 6720 1691 10560
rect -2229 6680 1691 6720
rect 2789 10560 6709 10600
rect 2789 6720 2829 10560
rect 6669 6720 6709 10560
rect 2789 6680 6709 6720
rect 7807 10560 11727 10600
rect 7807 6720 7847 10560
rect 11687 6720 11727 10560
rect 7807 6680 11727 6720
rect -12265 6240 -8345 6280
rect -12265 2400 -12225 6240
rect -8385 2400 -8345 6240
rect -12265 2360 -8345 2400
rect -7247 6240 -3327 6280
rect -7247 2400 -7207 6240
rect -3367 2400 -3327 6240
rect -7247 2360 -3327 2400
rect -2229 6240 1691 6280
rect -2229 2400 -2189 6240
rect 1651 2400 1691 6240
rect -2229 2360 1691 2400
rect 2789 6240 6709 6280
rect 2789 2400 2829 6240
rect 6669 2400 6709 6240
rect 2789 2360 6709 2400
rect 7807 6240 11727 6280
rect 7807 2400 7847 6240
rect 11687 2400 11727 6240
rect 7807 2360 11727 2400
rect -12265 1920 -8345 1960
rect -12265 -1920 -12225 1920
rect -8385 -1920 -8345 1920
rect -12265 -1960 -8345 -1920
rect -7247 1920 -3327 1960
rect -7247 -1920 -7207 1920
rect -3367 -1920 -3327 1920
rect -7247 -1960 -3327 -1920
rect -2229 1920 1691 1960
rect -2229 -1920 -2189 1920
rect 1651 -1920 1691 1920
rect -2229 -1960 1691 -1920
rect 2789 1920 6709 1960
rect 2789 -1920 2829 1920
rect 6669 -1920 6709 1920
rect 2789 -1960 6709 -1920
rect 7807 1920 11727 1960
rect 7807 -1920 7847 1920
rect 11687 -1920 11727 1920
rect 7807 -1960 11727 -1920
rect -12265 -2400 -8345 -2360
rect -12265 -6240 -12225 -2400
rect -8385 -6240 -8345 -2400
rect -12265 -6280 -8345 -6240
rect -7247 -2400 -3327 -2360
rect -7247 -6240 -7207 -2400
rect -3367 -6240 -3327 -2400
rect -7247 -6280 -3327 -6240
rect -2229 -2400 1691 -2360
rect -2229 -6240 -2189 -2400
rect 1651 -6240 1691 -2400
rect -2229 -6280 1691 -6240
rect 2789 -2400 6709 -2360
rect 2789 -6240 2829 -2400
rect 6669 -6240 6709 -2400
rect 2789 -6280 6709 -6240
rect 7807 -2400 11727 -2360
rect 7807 -6240 7847 -2400
rect 11687 -6240 11727 -2400
rect 7807 -6280 11727 -6240
rect -12265 -6720 -8345 -6680
rect -12265 -10560 -12225 -6720
rect -8385 -10560 -8345 -6720
rect -12265 -10600 -8345 -10560
rect -7247 -6720 -3327 -6680
rect -7247 -10560 -7207 -6720
rect -3367 -10560 -3327 -6720
rect -7247 -10600 -3327 -10560
rect -2229 -6720 1691 -6680
rect -2229 -10560 -2189 -6720
rect 1651 -10560 1691 -6720
rect -2229 -10600 1691 -10560
rect 2789 -6720 6709 -6680
rect 2789 -10560 2829 -6720
rect 6669 -10560 6709 -6720
rect 2789 -10600 6709 -10560
rect 7807 -6720 11727 -6680
rect 7807 -10560 7847 -6720
rect 11687 -10560 11727 -6720
rect 7807 -10600 11727 -10560
<< mimcap2contact >>
rect -12225 6720 -8385 10560
rect -7207 6720 -3367 10560
rect -2189 6720 1651 10560
rect 2829 6720 6669 10560
rect 7847 6720 11687 10560
rect -12225 2400 -8385 6240
rect -7207 2400 -3367 6240
rect -2189 2400 1651 6240
rect 2829 2400 6669 6240
rect 7847 2400 11687 6240
rect -12225 -1920 -8385 1920
rect -7207 -1920 -3367 1920
rect -2189 -1920 1651 1920
rect 2829 -1920 6669 1920
rect 7847 -1920 11687 1920
rect -12225 -6240 -8385 -2400
rect -7207 -6240 -3367 -2400
rect -2189 -6240 1651 -2400
rect 2829 -6240 6669 -2400
rect 7847 -6240 11687 -2400
rect -12225 -10560 -8385 -6720
rect -7207 -10560 -3367 -6720
rect -2189 -10560 1651 -6720
rect 2829 -10560 6669 -6720
rect 7847 -10560 11687 -6720
<< metal5 >>
rect -10465 10584 -10145 10800
rect -8025 10639 -7705 10800
rect -12249 10560 -8361 10584
rect -12249 6720 -12225 10560
rect -8385 6720 -8361 10560
rect -12249 6696 -8361 6720
rect -10465 6264 -10145 6696
rect -8025 6641 -7983 10639
rect -7747 6641 -7705 10639
rect -5447 10584 -5127 10800
rect -3007 10639 -2687 10800
rect -7231 10560 -3343 10584
rect -7231 6720 -7207 10560
rect -3367 6720 -3343 10560
rect -7231 6696 -3343 6720
rect -8025 6319 -7705 6641
rect -12249 6240 -8361 6264
rect -12249 2400 -12225 6240
rect -8385 2400 -8361 6240
rect -12249 2376 -8361 2400
rect -10465 1944 -10145 2376
rect -8025 2321 -7983 6319
rect -7747 2321 -7705 6319
rect -5447 6264 -5127 6696
rect -3007 6641 -2965 10639
rect -2729 6641 -2687 10639
rect -429 10584 -109 10800
rect 2011 10639 2331 10800
rect -2213 10560 1675 10584
rect -2213 6720 -2189 10560
rect 1651 6720 1675 10560
rect -2213 6696 1675 6720
rect -3007 6319 -2687 6641
rect -7231 6240 -3343 6264
rect -7231 2400 -7207 6240
rect -3367 2400 -3343 6240
rect -7231 2376 -3343 2400
rect -8025 1999 -7705 2321
rect -12249 1920 -8361 1944
rect -12249 -1920 -12225 1920
rect -8385 -1920 -8361 1920
rect -12249 -1944 -8361 -1920
rect -10465 -2376 -10145 -1944
rect -8025 -1999 -7983 1999
rect -7747 -1999 -7705 1999
rect -5447 1944 -5127 2376
rect -3007 2321 -2965 6319
rect -2729 2321 -2687 6319
rect -429 6264 -109 6696
rect 2011 6641 2053 10639
rect 2289 6641 2331 10639
rect 4589 10584 4909 10800
rect 7029 10639 7349 10800
rect 2805 10560 6693 10584
rect 2805 6720 2829 10560
rect 6669 6720 6693 10560
rect 2805 6696 6693 6720
rect 2011 6319 2331 6641
rect -2213 6240 1675 6264
rect -2213 2400 -2189 6240
rect 1651 2400 1675 6240
rect -2213 2376 1675 2400
rect -3007 1999 -2687 2321
rect -7231 1920 -3343 1944
rect -7231 -1920 -7207 1920
rect -3367 -1920 -3343 1920
rect -7231 -1944 -3343 -1920
rect -8025 -2321 -7705 -1999
rect -12249 -2400 -8361 -2376
rect -12249 -6240 -12225 -2400
rect -8385 -6240 -8361 -2400
rect -12249 -6264 -8361 -6240
rect -10465 -6696 -10145 -6264
rect -8025 -6319 -7983 -2321
rect -7747 -6319 -7705 -2321
rect -5447 -2376 -5127 -1944
rect -3007 -1999 -2965 1999
rect -2729 -1999 -2687 1999
rect -429 1944 -109 2376
rect 2011 2321 2053 6319
rect 2289 2321 2331 6319
rect 4589 6264 4909 6696
rect 7029 6641 7071 10639
rect 7307 6641 7349 10639
rect 9607 10584 9927 10800
rect 12047 10639 12367 10800
rect 7823 10560 11711 10584
rect 7823 6720 7847 10560
rect 11687 6720 11711 10560
rect 7823 6696 11711 6720
rect 7029 6319 7349 6641
rect 2805 6240 6693 6264
rect 2805 2400 2829 6240
rect 6669 2400 6693 6240
rect 2805 2376 6693 2400
rect 2011 1999 2331 2321
rect -2213 1920 1675 1944
rect -2213 -1920 -2189 1920
rect 1651 -1920 1675 1920
rect -2213 -1944 1675 -1920
rect -3007 -2321 -2687 -1999
rect -7231 -2400 -3343 -2376
rect -7231 -6240 -7207 -2400
rect -3367 -6240 -3343 -2400
rect -7231 -6264 -3343 -6240
rect -8025 -6641 -7705 -6319
rect -12249 -6720 -8361 -6696
rect -12249 -10560 -12225 -6720
rect -8385 -10560 -8361 -6720
rect -12249 -10584 -8361 -10560
rect -10465 -10800 -10145 -10584
rect -8025 -10639 -7983 -6641
rect -7747 -10639 -7705 -6641
rect -5447 -6696 -5127 -6264
rect -3007 -6319 -2965 -2321
rect -2729 -6319 -2687 -2321
rect -429 -2376 -109 -1944
rect 2011 -1999 2053 1999
rect 2289 -1999 2331 1999
rect 4589 1944 4909 2376
rect 7029 2321 7071 6319
rect 7307 2321 7349 6319
rect 9607 6264 9927 6696
rect 12047 6641 12089 10639
rect 12325 6641 12367 10639
rect 12047 6319 12367 6641
rect 7823 6240 11711 6264
rect 7823 2400 7847 6240
rect 11687 2400 11711 6240
rect 7823 2376 11711 2400
rect 7029 1999 7349 2321
rect 2805 1920 6693 1944
rect 2805 -1920 2829 1920
rect 6669 -1920 6693 1920
rect 2805 -1944 6693 -1920
rect 2011 -2321 2331 -1999
rect -2213 -2400 1675 -2376
rect -2213 -6240 -2189 -2400
rect 1651 -6240 1675 -2400
rect -2213 -6264 1675 -6240
rect -3007 -6641 -2687 -6319
rect -7231 -6720 -3343 -6696
rect -7231 -10560 -7207 -6720
rect -3367 -10560 -3343 -6720
rect -7231 -10584 -3343 -10560
rect -8025 -10800 -7705 -10639
rect -5447 -10800 -5127 -10584
rect -3007 -10639 -2965 -6641
rect -2729 -10639 -2687 -6641
rect -429 -6696 -109 -6264
rect 2011 -6319 2053 -2321
rect 2289 -6319 2331 -2321
rect 4589 -2376 4909 -1944
rect 7029 -1999 7071 1999
rect 7307 -1999 7349 1999
rect 9607 1944 9927 2376
rect 12047 2321 12089 6319
rect 12325 2321 12367 6319
rect 12047 1999 12367 2321
rect 7823 1920 11711 1944
rect 7823 -1920 7847 1920
rect 11687 -1920 11711 1920
rect 7823 -1944 11711 -1920
rect 7029 -2321 7349 -1999
rect 2805 -2400 6693 -2376
rect 2805 -6240 2829 -2400
rect 6669 -6240 6693 -2400
rect 2805 -6264 6693 -6240
rect 2011 -6641 2331 -6319
rect -2213 -6720 1675 -6696
rect -2213 -10560 -2189 -6720
rect 1651 -10560 1675 -6720
rect -2213 -10584 1675 -10560
rect -3007 -10800 -2687 -10639
rect -429 -10800 -109 -10584
rect 2011 -10639 2053 -6641
rect 2289 -10639 2331 -6641
rect 4589 -6696 4909 -6264
rect 7029 -6319 7071 -2321
rect 7307 -6319 7349 -2321
rect 9607 -2376 9927 -1944
rect 12047 -1999 12089 1999
rect 12325 -1999 12367 1999
rect 12047 -2321 12367 -1999
rect 7823 -2400 11711 -2376
rect 7823 -6240 7847 -2400
rect 11687 -6240 11711 -2400
rect 7823 -6264 11711 -6240
rect 7029 -6641 7349 -6319
rect 2805 -6720 6693 -6696
rect 2805 -10560 2829 -6720
rect 6669 -10560 6693 -6720
rect 2805 -10584 6693 -10560
rect 2011 -10800 2331 -10639
rect 4589 -10800 4909 -10584
rect 7029 -10639 7071 -6641
rect 7307 -10639 7349 -6641
rect 9607 -6696 9927 -6264
rect 12047 -6319 12089 -2321
rect 12325 -6319 12367 -2321
rect 12047 -6641 12367 -6319
rect 7823 -6720 11711 -6696
rect 7823 -10560 7847 -6720
rect 11687 -10560 11711 -6720
rect 7823 -10584 11711 -10560
rect 7029 -10800 7349 -10639
rect 9607 -10800 9927 -10584
rect 12047 -10639 12089 -6641
rect 12325 -10639 12367 -6641
rect 12047 -10800 12367 -10639
<< properties >>
string FIXED_BBOX 7727 6600 11807 10680
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 19.6 l 19.6 val 783.216 carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
