magic
tech sky130A
magscale 1 2
timestamp 1668729649
<< psubdiff >>
rect 8076 160 8100 370
rect 8380 160 8404 370
<< psubdiffcont >>
rect 8100 160 8380 370
<< locali >>
rect 7583 2169 7690 2211
rect 8084 160 8100 370
rect 8380 160 8396 370
<< viali >>
rect 5540 2160 5600 2200
rect 7280 2150 7340 2210
rect 7690 2160 7740 2220
rect 5840 2080 5892 2132
rect 8100 160 8380 370
<< metal1 >>
rect 6300 5000 6500 5400
rect 6620 5000 6820 5400
rect 6960 5000 7160 5400
rect 7580 5000 7780 5400
rect 7920 5020 8120 5420
rect 8240 5000 8440 5400
rect 4640 3300 6330 3500
rect 6440 3280 6640 3680
rect 6780 3260 6980 3660
rect 7100 3260 7640 3700
rect 8380 3690 8480 3700
rect 7760 3280 7960 3680
rect 8080 3280 8280 3680
rect 8380 3620 8400 3690
rect 8480 3620 8490 3690
rect 8380 3580 8480 3620
rect 8380 3510 8400 3580
rect 8480 3510 8490 3580
rect 8380 3470 8480 3510
rect 8380 3400 8390 3470
rect 8470 3400 8480 3470
rect 8380 3350 8480 3400
rect 8380 3280 8390 3350
rect 8470 3280 8480 3350
rect 7300 3060 7420 3260
rect 8680 3160 8920 3180
rect 8680 3060 8700 3160
rect 7300 2940 8700 3060
rect 4640 2820 4840 2860
rect 4640 2720 5640 2820
rect 4640 2660 4840 2720
rect 5540 2460 5640 2720
rect 8260 2660 8360 2940
rect 8680 2860 8700 2940
rect 8900 2860 8920 3160
rect 8680 2840 8920 2860
rect 8140 2600 8290 2610
rect 4640 2280 5260 2310
rect 4640 2160 4880 2280
rect 5010 2160 5090 2280
rect 5220 2160 5260 2280
rect 7680 2230 7790 2240
rect 4640 2120 5260 2160
rect 5360 2200 5620 2220
rect 5360 2160 5540 2200
rect 5600 2160 5620 2200
rect 5360 2140 5620 2160
rect 7268 2210 7352 2216
rect 7268 2150 7280 2210
rect 7340 2150 7352 2210
rect 7268 2144 7352 2150
rect 7680 2150 7690 2230
rect 7780 2150 7790 2230
rect 4640 2110 4840 2120
rect 5360 1610 5460 2140
rect 5830 2138 5840 2142
rect 5828 2130 5840 2138
rect 5892 2138 5902 2142
rect 7680 2140 7790 2150
rect 5820 2080 5840 2130
rect 5892 2130 5904 2138
rect 7000 2130 7060 2140
rect 5892 2080 5910 2130
rect 5828 2074 5904 2080
rect 7000 2060 7790 2110
rect 4640 1228 4840 1280
rect 5363 1228 5458 1610
rect 4640 1133 5458 1228
rect 4640 1080 4840 1133
rect 5640 60 5720 1980
rect 7700 60 7790 2060
rect 8130 2020 8290 2600
rect 8330 2020 8850 2600
rect 8130 1781 8180 2020
rect 8130 1780 8195 1781
rect 8110 1775 8220 1780
rect 8110 1685 8124 1775
rect 8214 1685 8220 1775
rect 8110 1680 8220 1685
rect 8130 1679 8195 1680
rect 8130 1400 8180 1679
rect 8260 1440 8360 1980
rect 8130 1210 8290 1400
rect 8340 1230 8530 1400
rect 8280 1120 8340 1180
rect 8430 860 8530 1230
rect 8140 700 8530 860
rect 8140 390 8310 700
rect 8060 370 8450 390
rect 8060 160 8100 370
rect 8380 160 8450 370
rect 8060 140 8450 160
rect 8140 60 8310 140
rect 8700 60 8850 2020
rect 5590 -140 5790 60
rect 7650 -140 7850 60
rect 8120 -140 8320 60
rect 8680 -140 8880 60
<< via1 >>
rect 8400 3620 8480 3690
rect 8400 3510 8480 3580
rect 8390 3400 8470 3470
rect 8390 3280 8470 3350
rect 8700 2860 8900 3160
rect 4880 2160 5010 2280
rect 5090 2160 5220 2280
rect 7280 2150 7340 2210
rect 7690 2220 7780 2230
rect 7690 2160 7740 2220
rect 7740 2160 7780 2220
rect 7690 2150 7780 2160
rect 5840 2132 5892 2142
rect 5840 2090 5892 2132
rect 8124 1685 8214 1775
<< metal2 >>
rect 7270 3810 8480 3890
rect 4840 2280 5260 2310
rect 4840 2160 4880 2280
rect 5010 2160 5090 2280
rect 5220 2160 5260 2280
rect 4840 2120 5260 2160
rect 7270 2210 7350 3810
rect 8400 3690 8480 3810
rect 8400 3580 8480 3620
rect 8400 3480 8480 3510
rect 8390 3470 8480 3480
rect 8470 3400 8480 3470
rect 8390 3390 8480 3400
rect 8400 3360 8480 3390
rect 8390 3350 8480 3360
rect 8470 3280 8480 3350
rect 8390 3270 8480 3280
rect 8680 3160 8920 3180
rect 8680 2860 8700 3160
rect 8900 2860 8920 3160
rect 8680 2840 8920 2860
rect 5840 2150 5892 2152
rect 7270 2150 7280 2210
rect 7340 2150 7350 2210
rect 5820 2142 5910 2150
rect 5820 2090 5840 2142
rect 5892 2090 5910 2142
rect 7270 2140 7350 2150
rect 7680 2230 7790 2240
rect 7680 2150 7690 2230
rect 7780 2150 7790 2230
rect 7680 2140 7790 2150
rect 5820 1775 5910 2090
rect 8110 1775 8220 1780
rect 5820 1685 8124 1775
rect 8214 1685 8220 1775
rect 8110 1680 8220 1685
<< via2 >>
rect 4880 2160 5010 2280
rect 5090 2160 5220 2280
rect 8700 2860 8900 3160
rect 7690 2150 7780 2230
<< metal3 >>
rect 8680 3160 8920 3180
rect 8680 2860 8700 3160
rect 8900 2860 8920 3160
rect 8680 2840 8920 2860
rect 4860 2280 5290 2300
rect 4860 2160 4880 2280
rect 5010 2160 5090 2280
rect 5220 2240 5290 2280
rect 5220 2230 7790 2240
rect 5220 2160 7690 2230
rect 4860 2150 7690 2160
rect 7780 2150 7790 2230
rect 4860 2140 7790 2150
rect 4860 2120 5290 2140
<< via3 >>
rect 8700 2860 8900 3160
<< metal4 >>
rect 8680 3160 9680 3180
rect 8680 2860 8700 3160
rect 8900 2860 9680 3160
rect 8680 2840 9680 2860
use sky130_fd_pr__cap_mim_m3_1_A4KLY5  XC1
timestamp 1667782711
transform 1 0 11770 0 1 3020
box -2870 -2820 2869 2820
use sky130_fd_pr__nfet_01v8_648S5X  XN1
timestamp 1667782711
transform 1 0 8311 0 1 1310
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGSNAL  XP1
timestamp 1667782711
transform 1 0 8311 0 1 2319
box -211 -519 211 519
use sky130_fd_pr__res_xhigh_po_0p35_RGJZ8N  XR2
timestamp 1667790215
transform 1 0 8016 0 1 4348
box -616 -1248 616 1248
use sky130_fd_pr__res_xhigh_po_0p35_RGJZ8N  sky130_fd_pr__res_xhigh_po_0p35_RGJZ8N_0
timestamp 1667790215
transform 1 0 6716 0 1 4348
box -616 -1248 616 1248
use sky130_fd_sc_hd__dfrbp_1  x1 ~/sky130_workspace-centos7/open_pdks/sky130/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5538 0 1 1948
box -38 -48 2154 592
<< labels >>
flabel metal1 4640 1080 4840 1280 0 FreeSans 256 0 0 0 clk
port 2 nsew
flabel metal1 7650 -140 7850 60 0 FreeSans 256 0 0 0 reset_b_dff
port 4 nsew
flabel metal1 8120 -140 8320 60 0 FreeSans 256 0 0 0 gnd
port 1 nsew
flabel metal1 8680 -140 8880 60 0 FreeSans 256 0 0 0 vd
port 7 nsew
flabel metal1 5590 -140 5790 60 0 FreeSans 256 0 0 0 gnd_d
port 6 nsew
flabel metal1 4640 2110 4840 2310 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 4640 2660 4840 2860 0 FreeSans 256 0 0 0 vpwr
port 5 nsew
flabel metal1 4640 3300 4840 3500 0 FreeSans 256 0 0 0 in
port 0 nsew
<< end >>
