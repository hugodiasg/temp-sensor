magic
tech sky130A
magscale 1 2
timestamp 1675895675
<< metal4 >>
rect -15145 13439 -9407 13480
rect -15145 8321 -9663 13439
rect -9427 8321 -9407 13439
rect -15145 8280 -9407 8321
rect -9007 13439 -3269 13480
rect -9007 8321 -3525 13439
rect -3289 8321 -3269 13439
rect -9007 8280 -3269 8321
rect -2869 13439 2869 13480
rect -2869 8321 2613 13439
rect 2849 8321 2869 13439
rect -2869 8280 2869 8321
rect 3269 13439 9007 13480
rect 3269 8321 8751 13439
rect 8987 8321 9007 13439
rect 3269 8280 9007 8321
rect 9407 13439 15145 13480
rect 9407 8321 14889 13439
rect 15125 8321 15145 13439
rect 9407 8280 15145 8321
rect -15145 7999 -9407 8040
rect -15145 2881 -9663 7999
rect -9427 2881 -9407 7999
rect -15145 2840 -9407 2881
rect -9007 7999 -3269 8040
rect -9007 2881 -3525 7999
rect -3289 2881 -3269 7999
rect -9007 2840 -3269 2881
rect -2869 7999 2869 8040
rect -2869 2881 2613 7999
rect 2849 2881 2869 7999
rect -2869 2840 2869 2881
rect 3269 7999 9007 8040
rect 3269 2881 8751 7999
rect 8987 2881 9007 7999
rect 3269 2840 9007 2881
rect 9407 7999 15145 8040
rect 9407 2881 14889 7999
rect 15125 2881 15145 7999
rect 9407 2840 15145 2881
rect -15145 2559 -9407 2600
rect -15145 -2559 -9663 2559
rect -9427 -2559 -9407 2559
rect -15145 -2600 -9407 -2559
rect -9007 2559 -3269 2600
rect -9007 -2559 -3525 2559
rect -3289 -2559 -3269 2559
rect -9007 -2600 -3269 -2559
rect -2869 2559 2869 2600
rect -2869 -2559 2613 2559
rect 2849 -2559 2869 2559
rect -2869 -2600 2869 -2559
rect 3269 2559 9007 2600
rect 3269 -2559 8751 2559
rect 8987 -2559 9007 2559
rect 3269 -2600 9007 -2559
rect 9407 2559 15145 2600
rect 9407 -2559 14889 2559
rect 15125 -2559 15145 2559
rect 9407 -2600 15145 -2559
rect -15145 -2881 -9407 -2840
rect -15145 -7999 -9663 -2881
rect -9427 -7999 -9407 -2881
rect -15145 -8040 -9407 -7999
rect -9007 -2881 -3269 -2840
rect -9007 -7999 -3525 -2881
rect -3289 -7999 -3269 -2881
rect -9007 -8040 -3269 -7999
rect -2869 -2881 2869 -2840
rect -2869 -7999 2613 -2881
rect 2849 -7999 2869 -2881
rect -2869 -8040 2869 -7999
rect 3269 -2881 9007 -2840
rect 3269 -7999 8751 -2881
rect 8987 -7999 9007 -2881
rect 3269 -8040 9007 -7999
rect 9407 -2881 15145 -2840
rect 9407 -7999 14889 -2881
rect 15125 -7999 15145 -2881
rect 9407 -8040 15145 -7999
rect -15145 -8321 -9407 -8280
rect -15145 -13439 -9663 -8321
rect -9427 -13439 -9407 -8321
rect -15145 -13480 -9407 -13439
rect -9007 -8321 -3269 -8280
rect -9007 -13439 -3525 -8321
rect -3289 -13439 -3269 -8321
rect -9007 -13480 -3269 -13439
rect -2869 -8321 2869 -8280
rect -2869 -13439 2613 -8321
rect 2849 -13439 2869 -8321
rect -2869 -13480 2869 -13439
rect 3269 -8321 9007 -8280
rect 3269 -13439 8751 -8321
rect 8987 -13439 9007 -8321
rect 3269 -13480 9007 -13439
rect 9407 -8321 15145 -8280
rect 9407 -13439 14889 -8321
rect 15125 -13439 15145 -8321
rect 9407 -13480 15145 -13439
<< via4 >>
rect -9663 8321 -9427 13439
rect -3525 8321 -3289 13439
rect 2613 8321 2849 13439
rect 8751 8321 8987 13439
rect 14889 8321 15125 13439
rect -9663 2881 -9427 7999
rect -3525 2881 -3289 7999
rect 2613 2881 2849 7999
rect 8751 2881 8987 7999
rect 14889 2881 15125 7999
rect -9663 -2559 -9427 2559
rect -3525 -2559 -3289 2559
rect 2613 -2559 2849 2559
rect 8751 -2559 8987 2559
rect 14889 -2559 15125 2559
rect -9663 -7999 -9427 -2881
rect -3525 -7999 -3289 -2881
rect 2613 -7999 2849 -2881
rect 8751 -7999 8987 -2881
rect 14889 -7999 15125 -2881
rect -9663 -13439 -9427 -8321
rect -3525 -13439 -3289 -8321
rect 2613 -13439 2849 -8321
rect 8751 -13439 8987 -8321
rect 14889 -13439 15125 -8321
<< mimcap2 >>
rect -15065 13360 -10025 13400
rect -15065 8400 -15025 13360
rect -10065 8400 -10025 13360
rect -15065 8360 -10025 8400
rect -8927 13360 -3887 13400
rect -8927 8400 -8887 13360
rect -3927 8400 -3887 13360
rect -8927 8360 -3887 8400
rect -2789 13360 2251 13400
rect -2789 8400 -2749 13360
rect 2211 8400 2251 13360
rect -2789 8360 2251 8400
rect 3349 13360 8389 13400
rect 3349 8400 3389 13360
rect 8349 8400 8389 13360
rect 3349 8360 8389 8400
rect 9487 13360 14527 13400
rect 9487 8400 9527 13360
rect 14487 8400 14527 13360
rect 9487 8360 14527 8400
rect -15065 7920 -10025 7960
rect -15065 2960 -15025 7920
rect -10065 2960 -10025 7920
rect -15065 2920 -10025 2960
rect -8927 7920 -3887 7960
rect -8927 2960 -8887 7920
rect -3927 2960 -3887 7920
rect -8927 2920 -3887 2960
rect -2789 7920 2251 7960
rect -2789 2960 -2749 7920
rect 2211 2960 2251 7920
rect -2789 2920 2251 2960
rect 3349 7920 8389 7960
rect 3349 2960 3389 7920
rect 8349 2960 8389 7920
rect 3349 2920 8389 2960
rect 9487 7920 14527 7960
rect 9487 2960 9527 7920
rect 14487 2960 14527 7920
rect 9487 2920 14527 2960
rect -15065 2480 -10025 2520
rect -15065 -2480 -15025 2480
rect -10065 -2480 -10025 2480
rect -15065 -2520 -10025 -2480
rect -8927 2480 -3887 2520
rect -8927 -2480 -8887 2480
rect -3927 -2480 -3887 2480
rect -8927 -2520 -3887 -2480
rect -2789 2480 2251 2520
rect -2789 -2480 -2749 2480
rect 2211 -2480 2251 2480
rect -2789 -2520 2251 -2480
rect 3349 2480 8389 2520
rect 3349 -2480 3389 2480
rect 8349 -2480 8389 2480
rect 3349 -2520 8389 -2480
rect 9487 2480 14527 2520
rect 9487 -2480 9527 2480
rect 14487 -2480 14527 2480
rect 9487 -2520 14527 -2480
rect -15065 -2960 -10025 -2920
rect -15065 -7920 -15025 -2960
rect -10065 -7920 -10025 -2960
rect -15065 -7960 -10025 -7920
rect -8927 -2960 -3887 -2920
rect -8927 -7920 -8887 -2960
rect -3927 -7920 -3887 -2960
rect -8927 -7960 -3887 -7920
rect -2789 -2960 2251 -2920
rect -2789 -7920 -2749 -2960
rect 2211 -7920 2251 -2960
rect -2789 -7960 2251 -7920
rect 3349 -2960 8389 -2920
rect 3349 -7920 3389 -2960
rect 8349 -7920 8389 -2960
rect 3349 -7960 8389 -7920
rect 9487 -2960 14527 -2920
rect 9487 -7920 9527 -2960
rect 14487 -7920 14527 -2960
rect 9487 -7960 14527 -7920
rect -15065 -8400 -10025 -8360
rect -15065 -13360 -15025 -8400
rect -10065 -13360 -10025 -8400
rect -15065 -13400 -10025 -13360
rect -8927 -8400 -3887 -8360
rect -8927 -13360 -8887 -8400
rect -3927 -13360 -3887 -8400
rect -8927 -13400 -3887 -13360
rect -2789 -8400 2251 -8360
rect -2789 -13360 -2749 -8400
rect 2211 -13360 2251 -8400
rect -2789 -13400 2251 -13360
rect 3349 -8400 8389 -8360
rect 3349 -13360 3389 -8400
rect 8349 -13360 8389 -8400
rect 3349 -13400 8389 -13360
rect 9487 -8400 14527 -8360
rect 9487 -13360 9527 -8400
rect 14487 -13360 14527 -8400
rect 9487 -13400 14527 -13360
<< mimcap2contact >>
rect -15025 8400 -10065 13360
rect -8887 8400 -3927 13360
rect -2749 8400 2211 13360
rect 3389 8400 8349 13360
rect 9527 8400 14487 13360
rect -15025 2960 -10065 7920
rect -8887 2960 -3927 7920
rect -2749 2960 2211 7920
rect 3389 2960 8349 7920
rect 9527 2960 14487 7920
rect -15025 -2480 -10065 2480
rect -8887 -2480 -3927 2480
rect -2749 -2480 2211 2480
rect 3389 -2480 8349 2480
rect 9527 -2480 14487 2480
rect -15025 -7920 -10065 -2960
rect -8887 -7920 -3927 -2960
rect -2749 -7920 2211 -2960
rect 3389 -7920 8349 -2960
rect 9527 -7920 14487 -2960
rect -15025 -13360 -10065 -8400
rect -8887 -13360 -3927 -8400
rect -2749 -13360 2211 -8400
rect 3389 -13360 8349 -8400
rect 9527 -13360 14487 -8400
<< metal5 >>
rect -12705 13384 -12385 13600
rect -9705 13439 -9385 13600
rect -15049 13360 -10041 13384
rect -15049 8400 -15025 13360
rect -10065 8400 -10041 13360
rect -15049 8376 -10041 8400
rect -12705 7944 -12385 8376
rect -9705 8321 -9663 13439
rect -9427 8321 -9385 13439
rect -6567 13384 -6247 13600
rect -3567 13439 -3247 13600
rect -8911 13360 -3903 13384
rect -8911 8400 -8887 13360
rect -3927 8400 -3903 13360
rect -8911 8376 -3903 8400
rect -9705 7999 -9385 8321
rect -15049 7920 -10041 7944
rect -15049 2960 -15025 7920
rect -10065 2960 -10041 7920
rect -15049 2936 -10041 2960
rect -12705 2504 -12385 2936
rect -9705 2881 -9663 7999
rect -9427 2881 -9385 7999
rect -6567 7944 -6247 8376
rect -3567 8321 -3525 13439
rect -3289 8321 -3247 13439
rect -429 13384 -109 13600
rect 2571 13439 2891 13600
rect -2773 13360 2235 13384
rect -2773 8400 -2749 13360
rect 2211 8400 2235 13360
rect -2773 8376 2235 8400
rect -3567 7999 -3247 8321
rect -8911 7920 -3903 7944
rect -8911 2960 -8887 7920
rect -3927 2960 -3903 7920
rect -8911 2936 -3903 2960
rect -9705 2559 -9385 2881
rect -15049 2480 -10041 2504
rect -15049 -2480 -15025 2480
rect -10065 -2480 -10041 2480
rect -15049 -2504 -10041 -2480
rect -12705 -2936 -12385 -2504
rect -9705 -2559 -9663 2559
rect -9427 -2559 -9385 2559
rect -6567 2504 -6247 2936
rect -3567 2881 -3525 7999
rect -3289 2881 -3247 7999
rect -429 7944 -109 8376
rect 2571 8321 2613 13439
rect 2849 8321 2891 13439
rect 5709 13384 6029 13600
rect 8709 13439 9029 13600
rect 3365 13360 8373 13384
rect 3365 8400 3389 13360
rect 8349 8400 8373 13360
rect 3365 8376 8373 8400
rect 2571 7999 2891 8321
rect -2773 7920 2235 7944
rect -2773 2960 -2749 7920
rect 2211 2960 2235 7920
rect -2773 2936 2235 2960
rect -3567 2559 -3247 2881
rect -8911 2480 -3903 2504
rect -8911 -2480 -8887 2480
rect -3927 -2480 -3903 2480
rect -8911 -2504 -3903 -2480
rect -9705 -2881 -9385 -2559
rect -15049 -2960 -10041 -2936
rect -15049 -7920 -15025 -2960
rect -10065 -7920 -10041 -2960
rect -15049 -7944 -10041 -7920
rect -12705 -8376 -12385 -7944
rect -9705 -7999 -9663 -2881
rect -9427 -7999 -9385 -2881
rect -6567 -2936 -6247 -2504
rect -3567 -2559 -3525 2559
rect -3289 -2559 -3247 2559
rect -429 2504 -109 2936
rect 2571 2881 2613 7999
rect 2849 2881 2891 7999
rect 5709 7944 6029 8376
rect 8709 8321 8751 13439
rect 8987 8321 9029 13439
rect 11847 13384 12167 13600
rect 14847 13439 15167 13600
rect 9503 13360 14511 13384
rect 9503 8400 9527 13360
rect 14487 8400 14511 13360
rect 9503 8376 14511 8400
rect 8709 7999 9029 8321
rect 3365 7920 8373 7944
rect 3365 2960 3389 7920
rect 8349 2960 8373 7920
rect 3365 2936 8373 2960
rect 2571 2559 2891 2881
rect -2773 2480 2235 2504
rect -2773 -2480 -2749 2480
rect 2211 -2480 2235 2480
rect -2773 -2504 2235 -2480
rect -3567 -2881 -3247 -2559
rect -8911 -2960 -3903 -2936
rect -8911 -7920 -8887 -2960
rect -3927 -7920 -3903 -2960
rect -8911 -7944 -3903 -7920
rect -9705 -8321 -9385 -7999
rect -15049 -8400 -10041 -8376
rect -15049 -13360 -15025 -8400
rect -10065 -13360 -10041 -8400
rect -15049 -13384 -10041 -13360
rect -12705 -13600 -12385 -13384
rect -9705 -13439 -9663 -8321
rect -9427 -13439 -9385 -8321
rect -6567 -8376 -6247 -7944
rect -3567 -7999 -3525 -2881
rect -3289 -7999 -3247 -2881
rect -429 -2936 -109 -2504
rect 2571 -2559 2613 2559
rect 2849 -2559 2891 2559
rect 5709 2504 6029 2936
rect 8709 2881 8751 7999
rect 8987 2881 9029 7999
rect 11847 7944 12167 8376
rect 14847 8321 14889 13439
rect 15125 8321 15167 13439
rect 14847 7999 15167 8321
rect 9503 7920 14511 7944
rect 9503 2960 9527 7920
rect 14487 2960 14511 7920
rect 9503 2936 14511 2960
rect 8709 2559 9029 2881
rect 3365 2480 8373 2504
rect 3365 -2480 3389 2480
rect 8349 -2480 8373 2480
rect 3365 -2504 8373 -2480
rect 2571 -2881 2891 -2559
rect -2773 -2960 2235 -2936
rect -2773 -7920 -2749 -2960
rect 2211 -7920 2235 -2960
rect -2773 -7944 2235 -7920
rect -3567 -8321 -3247 -7999
rect -8911 -8400 -3903 -8376
rect -8911 -13360 -8887 -8400
rect -3927 -13360 -3903 -8400
rect -8911 -13384 -3903 -13360
rect -9705 -13600 -9385 -13439
rect -6567 -13600 -6247 -13384
rect -3567 -13439 -3525 -8321
rect -3289 -13439 -3247 -8321
rect -429 -8376 -109 -7944
rect 2571 -7999 2613 -2881
rect 2849 -7999 2891 -2881
rect 5709 -2936 6029 -2504
rect 8709 -2559 8751 2559
rect 8987 -2559 9029 2559
rect 11847 2504 12167 2936
rect 14847 2881 14889 7999
rect 15125 2881 15167 7999
rect 14847 2559 15167 2881
rect 9503 2480 14511 2504
rect 9503 -2480 9527 2480
rect 14487 -2480 14511 2480
rect 9503 -2504 14511 -2480
rect 8709 -2881 9029 -2559
rect 3365 -2960 8373 -2936
rect 3365 -7920 3389 -2960
rect 8349 -7920 8373 -2960
rect 3365 -7944 8373 -7920
rect 2571 -8321 2891 -7999
rect -2773 -8400 2235 -8376
rect -2773 -13360 -2749 -8400
rect 2211 -13360 2235 -8400
rect -2773 -13384 2235 -13360
rect -3567 -13600 -3247 -13439
rect -429 -13600 -109 -13384
rect 2571 -13439 2613 -8321
rect 2849 -13439 2891 -8321
rect 5709 -8376 6029 -7944
rect 8709 -7999 8751 -2881
rect 8987 -7999 9029 -2881
rect 11847 -2936 12167 -2504
rect 14847 -2559 14889 2559
rect 15125 -2559 15167 2559
rect 14847 -2881 15167 -2559
rect 9503 -2960 14511 -2936
rect 9503 -7920 9527 -2960
rect 14487 -7920 14511 -2960
rect 9503 -7944 14511 -7920
rect 8709 -8321 9029 -7999
rect 3365 -8400 8373 -8376
rect 3365 -13360 3389 -8400
rect 8349 -13360 8373 -8400
rect 3365 -13384 8373 -13360
rect 2571 -13600 2891 -13439
rect 5709 -13600 6029 -13384
rect 8709 -13439 8751 -8321
rect 8987 -13439 9029 -8321
rect 11847 -8376 12167 -7944
rect 14847 -7999 14889 -2881
rect 15125 -7999 15167 -2881
rect 14847 -8321 15167 -7999
rect 9503 -8400 14511 -8376
rect 9503 -13360 9527 -8400
rect 14487 -13360 14511 -8400
rect 9503 -13384 14511 -13360
rect 8709 -13600 9029 -13439
rect 11847 -13600 12167 -13384
rect 14847 -13439 14889 -8321
rect 15125 -13439 15167 -8321
rect 14847 -13600 15167 -13439
<< properties >>
string FIXED_BBOX 9407 8280 14607 13480
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.2 l 25.2 val 1.289k carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
