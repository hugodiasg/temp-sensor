magic
tech sky130A
magscale 1 2
timestamp 1644948615
<< metal4 >>
rect -2579 7559 2579 7600
rect -2579 2641 2323 7559
rect 2559 2641 2579 7559
rect -2579 2600 2579 2641
rect -2579 2459 2579 2500
rect -2579 -2459 2323 2459
rect 2559 -2459 2579 2459
rect -2579 -2500 2579 -2459
rect -2579 -2641 2579 -2600
rect -2579 -7559 2323 -2641
rect 2559 -7559 2579 -2641
rect -2579 -7600 2579 -7559
<< via4 >>
rect 2323 2641 2559 7559
rect 2323 -2459 2559 2459
rect 2323 -7559 2559 -2641
<< mimcap2 >>
rect -2479 7460 2321 7500
rect -2479 2740 -1967 7460
rect 1809 2740 2321 7460
rect -2479 2700 2321 2740
rect -2479 2360 2321 2400
rect -2479 -2360 -1967 2360
rect 1809 -2360 2321 2360
rect -2479 -2400 2321 -2360
rect -2479 -2740 2321 -2700
rect -2479 -7460 -1967 -2740
rect 1809 -7460 2321 -2740
rect -2479 -7500 2321 -7460
<< mimcap2contact >>
rect -1967 2740 1809 7460
rect -1967 -2360 1809 2360
rect -1967 -7460 1809 -2740
<< metal5 >>
rect -239 7484 81 7650
rect 2281 7559 2601 7650
rect -1991 7460 1833 7484
rect -1991 2740 -1967 7460
rect 1809 2740 1833 7460
rect -1991 2716 1833 2740
rect -239 2384 81 2716
rect 2281 2641 2323 7559
rect 2559 2641 2601 7559
rect 2281 2459 2601 2641
rect -1991 2360 1833 2384
rect -1991 -2360 -1967 2360
rect 1809 -2360 1833 2360
rect -1991 -2384 1833 -2360
rect -239 -2716 81 -2384
rect 2281 -2459 2323 2459
rect 2559 -2459 2601 2459
rect 2281 -2641 2601 -2459
rect -1991 -2740 1833 -2716
rect -1991 -7460 -1967 -2740
rect 1809 -7460 1833 -2740
rect -1991 -7484 1833 -7460
rect -239 -7650 81 -7484
rect 2281 -7559 2323 -2641
rect 2559 -7559 2601 -2641
rect 2281 -7650 2601 -7559
<< properties >>
string FIXED_BBOX -2579 2600 2421 7600
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24 l 24 val 1.17k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
