magic
tech sky130A
magscale 1 2
timestamp 1701443238
<< metal1 >>
rect 6000 33780 7320 33820
rect 6000 33500 6940 33780
rect 7260 33500 7320 33780
rect 6000 33480 7320 33500
rect 6040 33140 6240 33480
rect -80 11320 1580 11460
rect 1760 11320 1780 11460
rect -80 11300 1780 11320
rect -320 10720 120 10920
rect 1550 6760 13100 6780
rect 1040 6560 1240 6760
rect 1550 6560 1560 6760
rect 1760 6560 12880 6760
rect 13080 6560 13100 6760
rect 1030 6400 1040 6560
rect 1220 6400 1240 6560
rect 1040 6380 1240 6400
rect 8750 5540 8760 5900
rect 8960 5540 8970 5900
rect 17310 5700 17320 5880
rect 17500 5700 17510 5880
rect 3490 5320 3500 5480
rect 4000 5320 4010 5480
rect 12020 5400 14480 5420
rect 12020 5240 12040 5400
rect 12200 5240 13720 5400
rect 13840 5240 14300 5400
rect 14440 5240 14480 5400
rect 12020 5220 14480 5240
rect 14310 4160 14320 4320
rect 14460 4160 14470 4320
rect 3810 3420 3950 3520
rect 4040 3360 4370 3560
rect 4040 2900 4380 3100
rect 4560 3080 5560 3100
rect 12030 3080 12040 3240
rect 12200 3080 12210 3240
rect 4560 2920 5380 3080
rect 5540 2920 5560 3080
rect 4560 2900 5560 2920
rect 5370 1960 5380 2120
rect 5540 1960 5550 2120
rect 4980 1800 5560 1820
rect 4980 1640 5000 1800
rect 5120 1640 5560 1800
rect 4980 1620 5560 1640
rect 12870 1580 12880 1780
rect 13080 1580 14020 1780
rect 14160 1580 14500 1780
rect 14330 1280 14340 1420
rect 14460 1280 14470 1420
rect 13080 1100 14500 1120
rect 13070 920 13080 1100
rect 13260 920 14500 1100
rect 14330 360 14340 540
rect 14460 360 14470 540
rect 190 40 200 160
rect 480 40 490 160
rect 15830 140 15990 160
rect 14770 0 14930 140
rect 14970 0 15130 140
rect 15230 120 15390 140
rect 15450 120 15610 140
rect 15630 120 15640 140
rect 15190 40 15640 120
rect 15230 0 15390 40
rect 15450 0 15610 40
rect 15630 20 15640 40
rect 15900 120 15990 140
rect 16250 120 16410 140
rect 16450 120 16610 140
rect 15900 40 16610 120
rect 15900 20 15990 40
rect 15650 0 15810 20
rect 16030 -20 16190 40
rect 16250 0 16410 40
rect 16450 0 16610 40
rect 16630 0 16950 140
rect 58 -1616 16098 -1596
rect 58 -1756 198 -1616
rect -62 -1916 198 -1756
rect 458 -1636 16098 -1616
rect 458 -1696 15678 -1636
rect 458 -1916 1058 -1696
rect -62 -1956 1058 -1916
rect 58 -1976 1058 -1956
rect 1218 -1876 15678 -1696
rect 15878 -1876 16098 -1636
rect 1218 -1976 16098 -1876
rect 58 -2036 16098 -1976
rect 4958 -2160 5158 -2156
rect 4358 -2196 4558 -2176
rect 4348 -2296 4358 -2196
rect 4558 -2296 4568 -2196
rect 4360 -2580 4560 -2296
rect 4950 -2300 4960 -2160
rect 5160 -2300 5170 -2160
rect 13078 -2176 13278 -2156
rect 14298 -2176 14498 -2156
rect 13078 -2276 13098 -2176
rect 13258 -2276 13278 -2176
rect 4958 -2576 5158 -2300
rect 13078 -2576 13278 -2276
rect 13698 -2196 13858 -2176
rect 13698 -2276 13718 -2196
rect 13838 -2276 13858 -2196
rect 13698 -2376 13858 -2276
rect 14008 -2296 14018 -2176
rect 14178 -2296 14188 -2176
rect 14298 -2276 14318 -2176
rect 14478 -2276 14498 -2176
rect 13658 -2576 13858 -2376
rect 14018 -2376 14178 -2296
rect 14298 -2376 14498 -2276
rect 14018 -2576 14218 -2376
rect 14278 -2576 14478 -2376
<< via1 >>
rect 6940 33500 7260 33780
rect 1580 11320 1760 11460
rect 1560 6560 1760 6760
rect 12880 6560 13080 6760
rect 1040 6400 1220 6560
rect 8760 5540 8960 5900
rect 17320 5700 17500 5880
rect 3500 5320 4000 5480
rect 12040 5240 12200 5400
rect 13720 5240 13840 5400
rect 14300 5240 14440 5400
rect 14320 4160 14460 4320
rect 4380 2900 4560 3100
rect 12040 3080 12200 3240
rect 5380 2920 5540 3080
rect 5380 1960 5540 2120
rect 5000 1640 5120 1800
rect 12880 1580 13080 1780
rect 14020 1580 14160 1780
rect 14340 1280 14460 1420
rect 13080 920 13260 1100
rect 14340 360 14460 540
rect 200 40 480 160
rect 15640 20 15900 140
rect 198 -1916 458 -1616
rect 1058 -1976 1218 -1696
rect 15678 -1876 15878 -1636
rect 4358 -2296 4558 -2196
rect 4960 -2300 5160 -2160
rect 13098 -2276 13258 -2176
rect 13718 -2276 13838 -2196
rect 14018 -2296 14178 -2176
rect 14318 -2276 14478 -2176
<< metal2 >>
rect 6940 33780 7260 33790
rect 6940 33490 7260 33500
rect 1560 11460 1780 11500
rect 1560 11320 1580 11460
rect 1760 11320 1780 11460
rect 1560 6760 1780 11320
rect 1040 6560 1220 6570
rect 1760 6560 1780 6760
rect 12880 6760 13100 6780
rect 13080 6560 13100 6760
rect 1560 6550 1760 6560
rect 1040 6390 1220 6400
rect 8760 5900 8960 5910
rect 8760 5530 8960 5540
rect 3500 5480 4000 5490
rect 3500 5310 4000 5320
rect 12020 5400 12220 5420
rect 12020 5240 12040 5400
rect 12200 5240 12220 5400
rect 12020 3240 12220 5240
rect 4360 3100 4560 3134
rect 4360 2900 4380 3100
rect 160 160 500 180
rect 160 40 200 160
rect 480 40 500 160
rect 160 -1384 500 40
rect 4360 -1384 4560 2900
rect 5360 3080 5560 3100
rect 5360 2920 5380 3080
rect 5540 2920 5560 3080
rect 12020 3080 12040 3240
rect 12200 3080 12220 3240
rect 12020 3060 12220 3080
rect 5360 2120 5560 2920
rect 5360 1960 5380 2120
rect 5540 1960 5560 2120
rect 5360 1940 5560 1960
rect 158 -1616 500 -1384
rect 158 -1916 198 -1616
rect 458 -1734 500 -1616
rect 4358 -1634 4560 -1384
rect 4980 1800 5140 1820
rect 4980 1640 5000 1800
rect 5120 1640 5140 1800
rect 1058 -1696 1218 -1686
rect 458 -1916 498 -1734
rect 158 -1956 498 -1916
rect 1058 -1986 1218 -1976
rect 4358 -2196 4558 -1634
rect 4980 -2150 5140 1640
rect 12880 1780 13100 6560
rect 17320 5880 17500 5890
rect 17320 5690 17500 5700
rect 13080 1580 13100 1780
rect 13700 5400 13860 5420
rect 13700 5240 13720 5400
rect 13840 5240 13860 5400
rect 12880 1570 13080 1580
rect 13080 1100 13280 1120
rect 13260 920 13280 1100
rect 13080 -1384 13280 920
rect 13700 -1384 13860 5240
rect 14280 5400 14460 5420
rect 14280 5240 14300 5400
rect 14440 5240 14460 5400
rect 14280 4320 14460 5240
rect 14280 4160 14320 4320
rect 14280 4140 14460 4160
rect 14020 1780 14160 1790
rect 14160 1580 14180 1780
rect 14020 -1384 14180 1580
rect 14300 1420 14500 1460
rect 14300 1280 14340 1420
rect 14460 1280 14500 1420
rect 14300 540 14500 1280
rect 14300 360 14340 540
rect 14460 360 14500 540
rect 14300 -1384 14500 360
rect 15600 140 15940 200
rect 15600 20 15640 140
rect 15900 20 15940 140
rect 15600 -1384 15940 20
rect 13078 -1620 13280 -1384
rect 13698 -1620 13860 -1384
rect 14018 -1620 14180 -1384
rect 14298 -1620 14500 -1384
rect 4358 -2306 4558 -2296
rect 4960 -2160 5160 -2150
rect 13078 -2176 13278 -1620
rect 13078 -2276 13098 -2176
rect 13258 -2276 13278 -2176
rect 13078 -2296 13278 -2276
rect 13698 -2196 13858 -1620
rect 13698 -2276 13718 -2196
rect 13838 -2276 13858 -2196
rect 13698 -2296 13858 -2276
rect 14018 -2176 14178 -1620
rect 14298 -2176 14498 -1620
rect 15598 -1630 15940 -1384
rect 15598 -1636 15938 -1630
rect 15598 -1876 15678 -1636
rect 15878 -1876 15938 -1636
rect 15598 -1956 15938 -1876
rect 14298 -2276 14318 -2176
rect 14478 -2276 14498 -2176
rect 14298 -2296 14498 -2276
rect 4960 -2310 5160 -2300
rect 14018 -2306 14178 -2296
<< via2 >>
rect 6940 33500 7260 33780
rect 1040 6400 1220 6560
rect 8760 5540 8960 5900
rect 3500 5320 4000 5480
rect 1058 -1976 1218 -1696
rect 17320 5700 17500 5880
<< metal3 >>
rect 6930 33780 7270 33785
rect 6930 33500 6940 33780
rect 7260 33500 7270 33780
rect 6930 33495 7270 33500
rect 1040 6565 1240 6580
rect 1030 6560 1240 6565
rect 1030 6400 1040 6560
rect 1220 6400 1240 6560
rect 1030 6395 1240 6400
rect 1040 -1384 1240 6395
rect 6980 5920 17520 5940
rect 6980 5720 7000 5920
rect 7260 5900 17520 5920
rect 7260 5720 8760 5900
rect 6980 5700 8760 5720
rect 8720 5540 8760 5700
rect 8960 5880 17520 5900
rect 8960 5700 17320 5880
rect 17500 5700 17520 5880
rect 8960 5540 9000 5700
rect 17310 5695 17510 5700
rect 8750 5535 8970 5540
rect 3490 5480 4010 5485
rect 3480 5320 3500 5480
rect 4000 5320 6920 5480
rect 3480 5300 6920 5320
rect 7240 5300 7250 5480
rect 3480 5280 7220 5300
rect 1038 -1634 1240 -1384
rect 1038 -1696 1238 -1634
rect 1038 -1976 1058 -1696
rect 1218 -1976 1238 -1696
rect 1038 -2036 1238 -1976
<< via3 >>
rect 6940 33500 7260 33780
rect 7000 5720 7260 5920
rect 6920 5300 7240 5480
<< metal4 >>
rect 6900 33780 7280 33860
rect 6900 33500 6940 33780
rect 7260 33500 7280 33780
rect 6900 6401 7280 33500
rect 6899 6279 7280 6401
rect 6900 5920 7280 6279
rect 6900 5720 7000 5920
rect 7260 5720 7280 5920
rect 6900 5480 7280 5720
rect 6900 5300 6920 5480
rect 7240 5300 7280 5480
rect 6900 5150 7280 5300
<< comment >>
rect 14280 -20 14300 0
use ask-modulator  ask-modulator_0 /foss/designs/temp-sensor/ask_modulator/mag
timestamp 1701402723
transform 1 0 -740 0 1 16920
box 660 -10360 31420 16420
use buffer  buffer_0 /foss/designs/temp-sensor/buffer/mag
timestamp 1700764089
transform 1 0 4468 0 1 -78
box 900 -1720 7760 5820
use sensor  sensor_0 /foss/designs/temp-sensor/sensor/mag
timestamp 1699935153
transform 1 0 660 0 1 2500
box -660 -2500 3580 3000
use sigma-delta  sigma-delta_0 /foss/designs/temp-sensor/sigma-delta_modulator/mag
timestamp 1701401593
transform 1 0 17480 0 1 520
box -3180 -520 12222 5680
<< labels >>
flabel metal1 6040 33620 6240 33820 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 -320 10720 -120 10920 0 FreeSans 1600 0 0 0 out
port 3 nsew
flabel metal1 4306 3508 4334 3538 0 FreeSans 1600 0 0 0 vtd
flabel metal1 11842 6654 11886 6698 0 FreeSans 800 0 0 0 out_sigma
flabel metal1 -62 -1956 138 -1756 0 FreeSans 1600 0 0 0 gnd
port 1 nsew
flabel metal1 14278 -2576 14478 -2376 0 FreeSans 1600 0 0 0 vpwr
port 4 nsew
flabel metal1 13078 -2576 13278 -2376 0 FreeSans 1600 0 0 0 clk
port 2 nsew
flabel metal1 13658 -2576 13858 -2376 0 FreeSans 1600 0 0 0 out_buff
port 7 nsew
flabel metal1 14018 -2576 14218 -2376 0 FreeSans 1600 0 0 0 out_sigma
port 9 nsew
flabel metal1 4958 -2576 5158 -2376 0 FreeSans 1600 0 0 0 ib
port 5 nsew
flabel metal1 4360 -2580 4560 -2380 0 FreeSans 1600 0 0 0 vts
port 8 nsew
<< end >>
