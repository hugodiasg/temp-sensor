magic
tech sky130A
magscale 1 2
timestamp 1657059275
<< nwell >>
rect -780 11500 -64 12434
rect -780 11160 -60 11500
rect 4900 11460 5616 12394
rect -780 10640 -64 11160
rect 4900 11120 5620 11460
rect 4900 10600 5616 11120
rect -780 9180 -64 10374
rect 460 9160 640 9380
<< pwell >>
rect -300 8360 356 9076
rect 5200 8200 6114 9616
<< mvnmos >>
rect -72 8618 128 8818
rect 5428 8458 5628 9358
rect 5686 8458 5886 9358
<< mvpmos >>
rect -522 10937 -322 12137
rect 5158 10897 5358 12097
rect -522 9477 -322 10077
<< mvndiff >>
rect -130 8806 -72 8818
rect -130 8630 -118 8806
rect -84 8630 -72 8806
rect -130 8618 -72 8630
rect 128 8806 186 8818
rect 128 8630 140 8806
rect 174 8630 186 8806
rect 128 8618 186 8630
rect 5370 9346 5428 9358
rect 5370 8470 5382 9346
rect 5416 8470 5428 9346
rect 5370 8458 5428 8470
rect 5628 9346 5686 9358
rect 5628 8470 5640 9346
rect 5674 8470 5686 9346
rect 5628 8458 5686 8470
rect 5886 9346 5944 9358
rect 5886 8470 5898 9346
rect 5932 8470 5944 9346
rect 5886 8458 5944 8470
<< mvpdiff >>
rect -580 12125 -522 12137
rect -580 10949 -568 12125
rect -534 10949 -522 12125
rect -580 10937 -522 10949
rect -322 12125 -264 12137
rect -322 10949 -310 12125
rect -276 10949 -264 12125
rect -322 10937 -264 10949
rect 5100 12085 5158 12097
rect 5100 10909 5112 12085
rect 5146 10909 5158 12085
rect 5100 10897 5158 10909
rect 5358 12085 5416 12097
rect 5358 10909 5370 12085
rect 5404 10909 5416 12085
rect 5358 10897 5416 10909
rect -580 10065 -522 10077
rect -580 9489 -568 10065
rect -534 9489 -522 10065
rect -580 9477 -522 9489
rect -322 10065 -264 10077
rect -322 9489 -310 10065
rect -276 9489 -264 10065
rect -322 9477 -264 9489
<< mvndiffc >>
rect -118 8630 -84 8806
rect 140 8630 174 8806
rect 5382 8470 5416 9346
rect 5640 8470 5674 9346
rect 5898 8470 5932 9346
<< mvpdiffc >>
rect -568 10949 -534 12125
rect -310 10949 -276 12125
rect 5112 10909 5146 12085
rect 5370 10909 5404 12085
rect -568 9489 -534 10065
rect -310 9489 -276 10065
<< mvpsubdiff >>
rect 5236 9568 6078 9580
rect 5236 9534 5344 9568
rect 5970 9534 6078 9568
rect 5236 9522 6078 9534
rect 5236 9472 5294 9522
rect -264 9028 320 9040
rect -264 8994 -156 9028
rect 212 8994 320 9028
rect -264 8982 320 8994
rect -264 8932 -206 8982
rect -264 8504 -252 8932
rect -218 8504 -206 8932
rect 262 8932 320 8982
rect -264 8454 -206 8504
rect 262 8504 274 8932
rect 308 8504 320 8932
rect 262 8454 320 8504
rect -264 8442 320 8454
rect -264 8408 -156 8442
rect 212 8408 320 8442
rect -264 8396 320 8408
rect 5236 8344 5248 9472
rect 5282 8344 5294 9472
rect 6020 9472 6078 9522
rect 5236 8294 5294 8344
rect 6020 8344 6032 9472
rect 6066 8344 6078 9472
rect 6020 8294 6078 8344
rect 5236 8282 6078 8294
rect 5236 8248 5344 8282
rect 5970 8248 6078 8282
rect 5236 8236 6078 8248
<< mvnsubdiff >>
rect -714 12356 -130 12368
rect -714 12322 -606 12356
rect -238 12322 -130 12356
rect -714 12310 -130 12322
rect -714 12260 -656 12310
rect -714 10814 -702 12260
rect -668 10814 -656 12260
rect -188 12260 -130 12310
rect -714 10764 -656 10814
rect -188 10814 -176 12260
rect -142 10814 -130 12260
rect -188 10764 -130 10814
rect -714 10752 -130 10764
rect -714 10718 -606 10752
rect -238 10718 -130 10752
rect -714 10706 -130 10718
rect 4966 12316 5550 12328
rect 4966 12282 5074 12316
rect 5442 12282 5550 12316
rect 4966 12270 5550 12282
rect 4966 12220 5024 12270
rect 4966 10774 4978 12220
rect 5012 10774 5024 12220
rect 5492 12220 5550 12270
rect 4966 10724 5024 10774
rect 5492 10774 5504 12220
rect 5538 10774 5550 12220
rect 5492 10724 5550 10774
rect 4966 10712 5550 10724
rect 4966 10678 5074 10712
rect 5442 10678 5550 10712
rect 4966 10666 5550 10678
rect -714 10296 -130 10308
rect -714 10262 -606 10296
rect -238 10262 -130 10296
rect -714 10250 -130 10262
rect -714 10200 -656 10250
rect -714 9354 -702 10200
rect -668 9354 -656 10200
rect -188 10200 -130 10250
rect -714 9304 -656 9354
rect -188 9354 -176 10200
rect -142 9354 -130 10200
rect -188 9304 -130 9354
rect -714 9292 -130 9304
rect -714 9258 -606 9292
rect -238 9258 -130 9292
rect -714 9246 -130 9258
<< mvpsubdiffcont >>
rect 5344 9534 5970 9568
rect -156 8994 212 9028
rect -252 8504 -218 8932
rect 274 8504 308 8932
rect -156 8408 212 8442
rect 5248 8344 5282 9472
rect 6032 8344 6066 9472
rect 5344 8248 5970 8282
<< mvnsubdiffcont >>
rect -606 12322 -238 12356
rect -702 10814 -668 12260
rect -176 10814 -142 12260
rect -606 10718 -238 10752
rect 5074 12282 5442 12316
rect 4978 10774 5012 12220
rect 5504 10774 5538 12220
rect 5074 10678 5442 10712
rect -606 10262 -238 10296
rect -702 9354 -668 10200
rect -176 9354 -142 10200
rect -606 9258 -238 9292
<< poly >>
rect -522 12218 -322 12234
rect -522 12184 -506 12218
rect -338 12184 -322 12218
rect -522 12137 -322 12184
rect -522 10890 -322 10937
rect -522 10856 -506 10890
rect -338 10856 -322 10890
rect -522 10840 -322 10856
rect 5158 12178 5358 12194
rect 5158 12144 5174 12178
rect 5342 12144 5358 12178
rect 5158 12097 5358 12144
rect 5158 10850 5358 10897
rect 5158 10816 5174 10850
rect 5342 10816 5358 10850
rect 5158 10800 5358 10816
rect -522 10158 -322 10174
rect -522 10124 -506 10158
rect -338 10124 -322 10158
rect -522 10077 -322 10124
rect -522 9430 -322 9477
rect -522 9396 -506 9430
rect -338 9396 -322 9430
rect -522 9380 -322 9396
rect -72 8890 128 8906
rect -72 8856 -56 8890
rect 112 8856 128 8890
rect -72 8818 128 8856
rect -72 8580 128 8618
rect -72 8546 -56 8580
rect 112 8546 128 8580
rect -72 8530 128 8546
rect 5428 9430 5628 9446
rect 5428 9396 5444 9430
rect 5612 9396 5628 9430
rect 5428 9358 5628 9396
rect 5686 9430 5886 9446
rect 5686 9396 5702 9430
rect 5870 9396 5886 9430
rect 5686 9358 5886 9396
rect 5428 8420 5628 8458
rect 5428 8386 5444 8420
rect 5612 8386 5628 8420
rect 5428 8370 5628 8386
rect 5686 8420 5886 8458
rect 5686 8386 5702 8420
rect 5870 8386 5886 8420
rect 5686 8370 5886 8386
<< polycont >>
rect -506 12184 -338 12218
rect -506 10856 -338 10890
rect 5174 12144 5342 12178
rect 5174 10816 5342 10850
rect -506 10124 -338 10158
rect -506 9396 -338 9430
rect -56 8856 112 8890
rect -56 8546 112 8580
rect 5444 9396 5612 9430
rect 5702 9396 5870 9430
rect 5444 8386 5612 8420
rect 5702 8386 5870 8420
<< locali >>
rect -702 12322 -606 12356
rect -238 12322 -142 12356
rect -702 12260 -668 12322
rect -176 12260 -142 12322
rect -522 12184 -506 12218
rect -338 12184 -322 12218
rect -568 12125 -534 12141
rect -568 10933 -534 10949
rect -310 12125 -276 12141
rect -310 10933 -276 10949
rect -522 10856 -506 10890
rect -338 10856 -322 10890
rect -702 10752 -668 10814
rect -176 10752 -142 10814
rect -702 10718 -606 10752
rect -238 10718 -142 10752
rect 4978 12282 5074 12316
rect 5442 12282 5538 12316
rect 4978 12220 5012 12282
rect 5504 12220 5538 12282
rect 5158 12144 5174 12178
rect 5342 12144 5358 12178
rect 5112 12085 5146 12101
rect 5112 10893 5146 10909
rect 5370 12085 5404 12101
rect 5370 10893 5404 10909
rect 5158 10816 5174 10850
rect 5342 10816 5358 10850
rect 4978 10712 5012 10774
rect 5504 10712 5538 10774
rect 4978 10678 5074 10712
rect 5442 10678 5538 10712
rect -702 10262 -606 10296
rect -238 10262 -142 10296
rect -702 10200 -668 10262
rect -176 10200 -142 10262
rect -522 10124 -506 10158
rect -338 10124 -322 10158
rect -568 10065 -534 10081
rect -568 9473 -534 9489
rect -310 10065 -276 10081
rect -310 9473 -276 9489
rect -522 9396 -506 9430
rect -338 9396 -322 9430
rect -702 9292 -668 9354
rect -176 9292 -142 9354
rect -702 9258 -606 9292
rect -238 9258 -142 9292
rect 5248 9534 5344 9568
rect 5970 9534 6066 9568
rect 5248 9472 5282 9534
rect -252 8994 -156 9028
rect 212 8994 308 9028
rect -252 8932 -218 8994
rect 274 8932 308 8994
rect -72 8856 -56 8890
rect 112 8856 128 8890
rect -118 8806 -84 8822
rect -118 8614 -84 8630
rect 140 8806 174 8822
rect 140 8614 174 8630
rect -72 8546 -56 8580
rect 112 8546 128 8580
rect -252 8442 -218 8504
rect 274 8442 308 8504
rect -252 8408 -156 8442
rect 212 8408 308 8442
rect 6032 9472 6066 9534
rect 5428 9396 5444 9430
rect 5612 9396 5628 9430
rect 5686 9396 5702 9430
rect 5870 9396 5886 9430
rect 5382 9346 5416 9362
rect 5382 8454 5416 8470
rect 5640 9346 5674 9362
rect 5640 8454 5674 8470
rect 5898 9346 5932 9362
rect 5898 8454 5932 8470
rect 5428 8386 5444 8420
rect 5612 8386 5628 8420
rect 5686 8386 5702 8420
rect 5870 8386 5886 8420
rect 5248 8282 5282 8344
rect 6032 8282 6066 8344
rect 5248 8248 5344 8282
rect 5970 8248 6066 8282
<< metal1 >>
rect 2460 12760 2660 12960
rect 700 12700 4140 12760
rect 700 12020 760 12700
rect 1680 12020 1740 12700
rect 2320 12380 2380 12700
rect 2320 12320 3460 12380
rect 4080 12000 4140 12700
rect -1040 11340 160 11420
rect -1040 11220 -840 11340
rect 100 10860 160 11340
rect 980 11100 1100 11120
rect 980 11020 1000 11100
rect 1080 11080 1100 11100
rect 1080 11020 1420 11080
rect 2620 11040 2680 11420
rect 3140 11040 3200 11420
rect 3500 11040 3620 11060
rect 980 11000 1100 11020
rect 2620 10980 3520 11040
rect 3500 10960 3520 10980
rect 3600 10960 3620 11040
rect 400 10860 460 10960
rect 3500 10940 3620 10960
rect 100 10800 4380 10860
rect -1040 10460 -840 10520
rect 4420 10460 4480 11000
rect 5460 10460 5880 10520
rect -1040 10380 1640 10460
rect -1040 10320 -840 10380
rect 700 10040 760 10260
rect 980 10080 1100 10100
rect 1440 10080 1640 10380
rect 4420 10400 5880 10460
rect 980 10040 1000 10080
rect 680 10000 1000 10040
rect 1080 10040 1100 10080
rect 1080 10000 1420 10040
rect 680 9980 1420 10000
rect 4420 9940 4480 10400
rect 5460 10320 5880 10400
rect 400 9540 520 9560
rect 400 9460 420 9540
rect 500 9460 520 9540
rect 400 9440 520 9460
rect 1000 9540 1120 9560
rect 1000 9460 1020 9540
rect 1100 9460 1120 9540
rect 2300 9540 3120 9600
rect 1000 9440 1120 9460
rect -1040 9200 -840 9280
rect 460 9200 640 9380
rect -1040 9140 640 9200
rect -1040 9080 -840 9140
rect 1040 8920 1100 9440
rect 1680 9140 1740 9520
rect 2300 9140 2360 9540
rect 2660 9380 2860 9540
rect 2940 9380 3120 9540
rect 1680 9080 2360 9140
rect 2460 9260 4180 9320
rect 620 8860 1520 8920
rect -1040 8360 -840 8420
rect 540 8360 600 8820
rect 860 8600 920 8860
rect 1680 8820 1740 9080
rect 1240 8360 1300 8820
rect 1540 8740 1740 8820
rect 1540 8720 1760 8740
rect 1640 8640 1660 8720
rect 1740 8640 1760 8720
rect 1640 8620 1760 8640
rect 2460 8360 2520 9260
rect 3480 8840 3660 8860
rect 3480 8800 3500 8840
rect 2880 8740 3500 8800
rect 3480 8720 3500 8740
rect 3640 8760 3660 8840
rect 4180 8760 4380 8800
rect 3640 8720 4380 8760
rect 3480 8700 4380 8720
rect -1040 8300 2520 8360
rect -1040 8220 -840 8300
rect 2460 8240 2580 8300
<< via1 >>
rect 1000 11020 1080 11100
rect 3520 10960 3600 11040
rect 1000 10000 1080 10080
rect 420 9460 500 9540
rect 1020 9460 1100 9540
rect 1660 8640 1740 8720
rect 3500 8720 3640 8840
<< metal2 >>
rect 980 11100 1100 11120
rect 980 11020 1000 11100
rect 1080 11020 1100 11100
rect 980 11000 1100 11020
rect 3500 11040 3620 11060
rect 1000 10100 1060 11000
rect 3500 10960 3520 11040
rect 3600 10960 3620 11040
rect 3500 10940 3620 10960
rect 980 10080 1100 10100
rect 980 10000 1000 10080
rect 1080 10000 1100 10080
rect 980 9980 1100 10000
rect 400 9540 520 9560
rect 400 9460 420 9540
rect 500 9520 520 9540
rect 1000 9540 1120 9560
rect 1000 9520 1020 9540
rect 500 9460 1020 9520
rect 1100 9460 1120 9540
rect 400 9440 520 9460
rect 1000 9440 1120 9460
rect 3520 8860 3580 10940
rect 3480 8840 3660 8860
rect 1640 8720 1760 8740
rect 1640 8640 1660 8720
rect 1740 8640 1760 8720
rect 3480 8720 3500 8840
rect 3640 8720 3660 8840
rect 3480 8700 3660 8720
rect 1640 8620 1760 8640
rect 1660 8140 1720 8620
rect 1600 8120 1800 8140
rect 1600 8020 1620 8120
rect 1780 8020 1800 8120
rect 1600 8000 1800 8020
<< via2 >>
rect 3500 8720 3640 8840
rect 1620 8020 1780 8120
<< metal3 >>
rect 3480 8840 3660 8860
rect 3480 8720 3500 8840
rect 3640 8720 3660 8840
rect 3480 8700 3660 8720
rect 1600 8120 1800 8140
rect 1600 8020 1620 8120
rect 1780 8020 1800 8120
rect 1600 7660 1800 8020
<< via3 >>
rect 3500 8720 3640 8840
<< metal4 >>
rect 3480 8840 3660 8860
rect 3480 8720 3500 8840
rect 3640 8720 3660 8840
rect 3480 7680 3660 8720
use sky130_fd_pr__cap_mim_m3_1_2NYK3R  XCC
timestamp 1656875000
transform 1 0 2450 0 1 5800
box -2250 -2200 2249 2200
use sky130_fd_pr__pfet_g5v0d10v5_GYM5UZ  XM1
timestamp 1656875158
transform 1 0 558 0 1 9737
box -358 -597 358 597
use sky130_fd_pr__pfet_g5v0d10v5_G8J5UZ  XM2
timestamp 1656875158
transform 1 0 1538 0 1 9737
box -358 -597 358 597
use sky130_fd_pr__nfet_g5v0d10v5_9YTB7P  XM3
timestamp 1656875158
transform 1 0 728 0 1 8718
box -328 -358 328 358
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  XM5
timestamp 1656875000
transform 1 0 558 0 1 11497
box -358 -897 358 897
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  XM6
timestamp 1656875000
transform 1 0 1538 0 1 11497
box -358 -897 358 897
use sky130_fd_pr__nfet_g5v0d10v5_G8BGHZ  XM7
timestamp 1656875210
transform 1 0 2897 0 1 8908
box -457 -708 457 708
use sky130_fd_pr__pfet_g5v0d10v5_8C84A7  XM8
timestamp 1656875000
transform 1 0 2905 0 1 11647
box -745 -1047 745 1047
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  XM10
timestamp 1656875000
transform 1 0 4278 0 1 11497
box -358 -897 358 897
use sky130_fd_pr__nfet_g5v0d10v5_9YTB7P  sky130_fd_pr__nfet_g5v0d10v5_9YTB7P_0
timestamp 1656875158
transform 1 0 1428 0 1 8718
box -328 -358 328 358
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  sky130_fd_pr__pfet_g5v0d10v5_GYMD5T_0
timestamp 1656875000
transform 1 0 4278 0 1 9437
box -358 -897 358 897
<< labels >>
flabel metal1 2460 12760 2660 12960 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel space 1020 10580 1160 10620 0 FreeSans 800 0 0 0 b
flabel metal1 1080 9360 1080 9360 0 FreeSans 800 0 0 0 c
flabel metal2 1680 8220 1680 8220 0 FreeSans 800 0 0 0 d
flabel metal1 3400 8760 3400 8760 0 FreeSans 800 0 0 0 e
flabel metal1 -1040 11220 -840 11420 0 FreeSans 1600 0 0 0 ib
port 1 nsew
flabel metal1 -1040 8220 -840 8420 0 FreeSans 1600 0 0 0 vs
port 5 nsew
flabel metal1 -1040 9080 -840 9280 0 FreeSans 1600 0 0 0 in1
port 4 nsew
flabel metal1 -1040 10320 -840 10520 0 FreeSans 1600 0 0 0 in2
port 3 nsew
flabel metal1 5680 10320 5880 10520 0 FreeSans 1600 0 0 0 out
port 2 nsew
<< end >>
