magic
tech sky130A
magscale 1 2
timestamp 1700063261
<< nmos >>
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
<< ndiff >>
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
<< ndiffc >>
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
<< poly >>
rect -487 172 -287 188
rect -487 138 -471 172
rect -303 138 -287 172
rect -487 100 -287 138
rect -229 172 -29 188
rect -229 138 -213 172
rect -45 138 -29 172
rect -229 100 -29 138
rect 29 172 229 188
rect 29 138 45 172
rect 213 138 229 172
rect 29 100 229 138
rect 287 172 487 188
rect 287 138 303 172
rect 471 138 487 172
rect 287 100 487 138
rect -487 -138 -287 -100
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -487 -188 -287 -172
rect -229 -138 -29 -100
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect -229 -188 -29 -172
rect 29 -138 229 -100
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 29 -188 229 -172
rect 287 -138 487 -100
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 287 -188 487 -172
<< polycont >>
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
<< locali >>
rect -487 138 -471 172
rect -303 138 -287 172
rect -229 138 -213 172
rect -45 138 -29 172
rect 29 138 45 172
rect 213 138 229 172
rect 287 138 303 172
rect 471 138 487 172
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 287 -172 303 -138
rect 471 -172 487 -138
<< viali >>
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
<< metal1 >>
rect -483 172 -291 178
rect -483 138 -471 172
rect -303 138 -291 172
rect -483 132 -291 138
rect -225 172 -33 178
rect -225 138 -213 172
rect -45 138 -33 172
rect -225 132 -33 138
rect 33 172 225 178
rect 33 138 45 172
rect 213 138 225 172
rect 33 132 225 138
rect 291 172 483 178
rect 291 138 303 172
rect 471 138 483 172
rect 291 132 483 138
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect -483 -138 -291 -132
rect -483 -172 -471 -138
rect -303 -172 -291 -138
rect -483 -178 -291 -172
rect -225 -138 -33 -132
rect -225 -172 -213 -138
rect -45 -172 -33 -138
rect -225 -178 -33 -172
rect 33 -138 225 -132
rect 33 -172 45 -138
rect 213 -172 225 -138
rect 33 -178 225 -172
rect 291 -138 483 -132
rect 291 -172 303 -138
rect 471 -172 483 -138
rect 291 -178 483 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
