magic
tech sky130A
timestamp 1645034384
<< metal4 >>
rect -600 900 1500 1500
<< metal5 >>
rect 0 14400 15000 15000
rect 0 13500 14100 14100
rect 0 600 600 13500
rect 13500 1500 14100 13500
rect 900 900 14100 1500
rect 14400 600 15000 14400
rect 0 0 15000 600
<< end >>
