magic
tech sky130A
magscale 1 2
timestamp 1645556896
<< metal1 >>
rect 6340 -1740 9360 -1640
rect 6340 -2100 6380 -1740
rect 7100 -2100 9360 -1740
rect 6340 -2180 9360 -2100
rect 10360 -1720 12600 -1620
rect 10360 -2080 11840 -1720
rect 12560 -2080 12600 -1720
rect 10360 -2160 12600 -2080
rect 8480 -2800 8680 -2180
rect 8860 -2580 10360 -2240
rect 9960 -2800 10360 -2580
rect 6340 -4480 9760 -2800
rect 9880 -3360 10360 -2800
rect 9880 -3740 10660 -3360
rect 9880 -4480 10360 -3740
rect 9718 -4646 9884 -4572
rect 9720 -5160 9880 -4646
rect 6340 -5360 9880 -5160
rect 10480 -5980 10660 -3740
rect 6340 -6180 10660 -5980
rect 10960 -8520 11560 -2160
rect 6340 -9140 11560 -8520
<< via1 >>
rect 6380 -2100 7100 -1740
rect 11840 -2080 12560 -1720
<< metal2 >>
rect 6340 -1740 7140 -1700
rect 6340 -2100 6380 -1740
rect 7100 -2100 7140 -1740
rect 6340 -2180 7140 -2100
rect 11800 -1720 12600 -1680
rect 11800 -2080 11840 -1720
rect 12560 -2080 12600 -1720
rect 11800 -2160 12600 -2080
<< via2 >>
rect 6380 -2100 7100 -1740
rect 11840 -2080 12560 -1720
<< metal3 >>
rect 6340 -1740 7140 -1700
rect 6340 -2100 6380 -1740
rect 7100 -2100 7140 -1740
rect 6340 -2180 7140 -2100
rect 11800 -1720 12600 -1680
rect 11800 -2080 11840 -1720
rect 12560 -2080 12600 -1720
rect 11800 -2160 12600 -2080
<< via3 >>
rect 6380 -2100 7100 -1740
rect 11840 -2080 12560 -1720
<< metal4 >>
rect 6339 14620 11480 15820
rect 11660 14620 13744 15820
rect 6340 -1740 7140 14620
rect 9440 13538 10420 14620
rect 6340 -2100 6380 -1740
rect 7100 -2100 7140 -1740
rect 6340 -2180 7140 -2100
rect 11800 -1720 12600 -1680
rect 11800 -2080 11840 -1720
rect 12560 -2080 12600 -1720
rect 11800 -2160 12600 -2080
<< rmetal4 >>
rect 11480 14620 11660 15820
<< via4 >>
rect 11840 -2080 12560 -1720
<< metal5 >>
rect 9500 390 10300 400
rect 9500 -624 10336 390
rect 9500 -1034 10320 -624
rect 9500 -1060 12590 -1034
rect 9500 -1540 12600 -1060
rect 11800 -1720 12600 -1540
rect 11800 -2080 11840 -1720
rect 12560 -2080 12600 -1720
rect 11800 -11160 12600 -2080
rect 11800 -11180 12628 -11160
rect 11800 -12380 14944 -11180
use 1  1_0
timestamp 1645556896
transform 1 0 13744 0 -1 17620
box -1200 0 30000 30000
use sky130_fd_pr__cap_mim_m3_2_9XH3MC  sky130_fd_pr__cap_mim_m3_2_9XH3MC_0
timestamp 1645036902
transform -1 0 9984 0 1 6691
box -2514 -7455 2536 7455
use sky130_fd_pr__nfet_g5v0d10v5_PWYS4E  sky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0
timestamp 1644948032
transform 1 0 9796 0 1 -3646
box -278 -1128 278 1128
use sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN  sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0
timestamp 1644948032
transform 0 1 9872 -1 0 -2093
box -201 -1098 201 1098
<< labels >>
flabel metal1 6340 -6180 6540 -5980 0 FreeSans 128 0 0 0 gnd
port 0 nsew
flabel metal1 6340 -5360 6540 -5160 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 6340 -3040 6540 -2840 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 6340 -8720 6540 -8520 0 FreeSans 128 0 0 0 vd
port 3 nsew
<< end >>
