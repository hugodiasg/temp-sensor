magic
tech sky130A
magscale 1 2
timestamp 1645793055
<< metal4 >>
rect -2179 6359 2179 6400
rect -2179 2241 1923 6359
rect 2159 2241 2179 6359
rect -2179 2200 2179 2241
rect -2179 2059 2179 2100
rect -2179 -2059 1923 2059
rect 2159 -2059 2179 2059
rect -2179 -2100 2179 -2059
rect -2179 -2241 2179 -2200
rect -2179 -6359 1923 -2241
rect 2159 -6359 2179 -2241
rect -2179 -6400 2179 -6359
<< via4 >>
rect 1923 2241 2159 6359
rect 1923 -2059 2159 2059
rect 1923 -6359 2159 -2241
<< mimcap2 >>
rect -2079 6260 1921 6300
rect -2079 2340 -1647 6260
rect 1489 2340 1921 6260
rect -2079 2300 1921 2340
rect -2079 1960 1921 2000
rect -2079 -1960 -1647 1960
rect 1489 -1960 1921 1960
rect -2079 -2000 1921 -1960
rect -2079 -2340 1921 -2300
rect -2079 -6260 -1647 -2340
rect 1489 -6260 1921 -2340
rect -2079 -6300 1921 -6260
<< mimcap2contact >>
rect -1647 2340 1489 6260
rect -1647 -1960 1489 1960
rect -1647 -6260 1489 -2340
<< metal5 >>
rect -239 6284 81 6450
rect 1881 6359 2201 6450
rect -1671 6260 1513 6284
rect -1671 2340 -1647 6260
rect 1489 2340 1513 6260
rect -1671 2316 1513 2340
rect -239 1984 81 2316
rect 1881 2241 1923 6359
rect 2159 2241 2201 6359
rect 1881 2059 2201 2241
rect -1671 1960 1513 1984
rect -1671 -1960 -1647 1960
rect 1489 -1960 1513 1960
rect -1671 -1984 1513 -1960
rect -239 -2316 81 -1984
rect 1881 -2059 1923 2059
rect 2159 -2059 2201 2059
rect 1881 -2241 2201 -2059
rect -1671 -2340 1513 -2316
rect -1671 -6260 -1647 -2340
rect 1489 -6260 1513 -2340
rect -1671 -6284 1513 -6260
rect -239 -6450 81 -6284
rect 1881 -6359 1923 -2241
rect 2159 -6359 2201 -2241
rect 1881 -6450 2201 -6359
<< properties >>
string FIXED_BBOX -2179 2200 2021 6400
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
