magic
tech sky130A
magscale 1 2
timestamp 1646429306
<< mvpsubdiff >>
rect 406200 555400 408200 555424
rect 406200 552976 408200 553000
<< mvpsubdiffcont >>
rect 406200 553000 408200 555400
<< locali >>
rect 406200 555400 408200 555416
rect 406200 552984 408200 553000
<< viali >>
rect 406200 553000 408200 555400
<< metal1 >>
rect 404800 576600 417600 576800
rect 404800 575200 411200 576600
rect 417600 575200 417610 576600
rect 404800 575000 417600 575200
rect 404800 557800 413600 558000
rect 404800 555800 410400 557800
rect 413400 555800 413600 557800
rect 404800 555600 413600 555800
rect 406000 555400 408400 555600
rect 406000 553000 406200 555400
rect 408200 553000 408400 555400
rect 406000 552800 408400 553000
rect 404800 531400 412600 531600
rect 404800 529200 409800 531400
rect 412400 529200 412600 531400
rect 404800 529000 412600 529200
<< via1 >>
rect 411200 575200 417600 576600
rect 410400 555800 413400 557800
rect 409800 529200 412400 531400
<< metal2 >>
rect 411000 576600 417800 576800
rect 411000 575200 411200 576600
rect 417600 575200 417800 576600
rect 411000 575000 417800 575200
rect 408000 557800 413600 558000
rect 408000 555800 410400 557800
rect 413400 555800 413600 557800
rect 408000 555600 413600 555800
rect 409600 531400 412600 531600
rect 409600 529200 409800 531400
rect 412400 529200 412600 531400
rect 409600 529000 412600 529200
<< via2 >>
rect 411200 575200 417600 576600
rect 410400 555800 413400 557800
rect 409800 529200 412400 531400
<< metal3 >>
rect 411000 576600 417800 576800
rect 411000 575200 411200 576600
rect 417600 575200 417800 576600
rect 411000 575000 417800 575200
rect 408000 557800 413600 558000
rect 408000 555800 410400 557800
rect 413400 555800 413600 557800
rect 408000 555600 413600 555800
rect 409600 531400 412600 531600
rect 409600 529200 409800 531400
rect 412400 529200 412600 531400
rect 409600 529000 412600 529200
<< via3 >>
rect 411200 575200 417600 576600
rect 410400 555800 413400 557800
rect 409800 529200 412400 531400
<< metal4 >>
rect 411000 576600 417800 576800
rect 411000 575200 411200 576600
rect 417600 575200 417800 576600
rect 411000 575000 417800 575200
rect 415600 558000 418600 562200
rect 421200 558000 424200 562200
rect 426600 558000 429600 562200
rect 408000 557800 429600 558000
rect 408000 555800 410400 557800
rect 413400 555800 429600 557800
rect 448160 558780 449820 558800
rect 448160 557240 448180 558780
rect 449800 557240 449820 558780
rect 448160 557220 449820 557240
rect 408000 555600 429600 555800
rect 410200 552600 413200 555600
rect 415600 552000 418600 555600
rect 421200 551800 424200 555600
rect 426600 552400 429600 555600
rect 409600 531400 412600 531600
rect 409600 529200 409800 531400
rect 412400 529200 412600 531400
rect 409600 529000 412600 529200
<< via4 >>
rect 411200 575200 417600 576600
rect 448180 557240 449800 558780
rect 409800 529200 412400 531400
<< metal5 >>
rect 411000 576600 433250 576800
rect 411000 575200 411200 576600
rect 417600 575200 433250 576600
rect 411000 575000 433250 575200
rect 415975 574975 433250 575000
rect 415975 573175 417625 574975
rect 421600 573200 423250 574975
rect 427200 573200 428850 574975
rect 431600 571500 433250 574975
rect 431600 571180 433220 571200
rect 433240 571180 433250 571190
rect 431600 563200 433250 571180
rect 448168 558804 449820 558820
rect 448156 558780 449824 558804
rect 448156 557240 448180 558780
rect 449800 557240 449824 558780
rect 448156 557216 449824 557240
rect 410400 533425 412800 536000
rect 415600 533425 418600 536000
rect 421400 533425 424400 536000
rect 427000 533425 430000 536400
rect 448168 533800 449818 557216
rect 448168 533425 449800 533800
rect 410400 531800 449800 533425
rect 410400 531600 412600 531800
rect 436400 531775 447400 531800
rect 409600 531400 412600 531600
rect 409600 529200 409800 531400
rect 412400 529200 412600 531400
rect 409600 529000 412600 529200
<< rm5 >>
rect 431600 571200 433250 571500
rect 433220 571190 433250 571200
rect 433220 571180 433240 571190
use l0  l0_0
timestamp 1646185352
transform 1 0 388400 0 1 505600
box 43200 43200 60788 59200
use sky130_fd_pr__cap_mim_m3_2_4GE4YE  sky130_fd_pr__cap_mim_m3_2_4GE4YE_0
timestamp 1646428335
transform 1 0 416672 0 1 566721
box -2472 -7329 2494 7329
use sky130_fd_pr__cap_mim_m3_2_4GE4YE  sky130_fd_pr__cap_mim_m3_2_4GE4YE_1
timestamp 1646428335
transform 1 0 422472 0 1 566721
box -2472 -7329 2494 7329
use sky130_fd_pr__cap_mim_m3_2_4GE4YE  sky130_fd_pr__cap_mim_m3_2_4GE4YE_2
timestamp 1646428335
transform 1 0 428272 0 1 566721
box -2472 -7329 2494 7329
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_0
timestamp 1646428335
transform 1 0 411186 0 1 544626
box -2586 -10228 2608 10228
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_1
timestamp 1646428335
transform 1 0 416786 0 1 544626
box -2586 -10228 2608 10228
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_2
timestamp 1646428335
transform 1 0 422786 0 1 544626
box -2586 -10228 2608 10228
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_3
timestamp 1646428335
transform 1 0 428586 0 1 544626
box -2586 -10228 2608 10228
<< labels >>
flabel metal1 404800 529000 407200 531600 0 FreeSans 1600 0 0 0 out
port 4 nsew
flabel metal1 404800 575000 406600 576800 0 FreeSans 1600 0 0 0 in
port 5 nsew
flabel metal1 404800 556000 406600 557800 0 FreeSans 1600 0 0 0 gnd
port 2 nsew
<< end >>
