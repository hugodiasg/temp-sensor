magic
tech sky130A
magscale 1 2
timestamp 1675895675
<< metal4 >>
rect -14145 12439 -8807 12480
rect -14145 7721 -9063 12439
rect -8827 7721 -8807 12439
rect -14145 7680 -8807 7721
rect -8407 12439 -3069 12480
rect -8407 7721 -3325 12439
rect -3089 7721 -3069 12439
rect -8407 7680 -3069 7721
rect -2669 12439 2669 12480
rect -2669 7721 2413 12439
rect 2649 7721 2669 12439
rect -2669 7680 2669 7721
rect 3069 12439 8407 12480
rect 3069 7721 8151 12439
rect 8387 7721 8407 12439
rect 3069 7680 8407 7721
rect 8807 12439 14145 12480
rect 8807 7721 13889 12439
rect 14125 7721 14145 12439
rect 8807 7680 14145 7721
rect -14145 7399 -8807 7440
rect -14145 2681 -9063 7399
rect -8827 2681 -8807 7399
rect -14145 2640 -8807 2681
rect -8407 7399 -3069 7440
rect -8407 2681 -3325 7399
rect -3089 2681 -3069 7399
rect -8407 2640 -3069 2681
rect -2669 7399 2669 7440
rect -2669 2681 2413 7399
rect 2649 2681 2669 7399
rect -2669 2640 2669 2681
rect 3069 7399 8407 7440
rect 3069 2681 8151 7399
rect 8387 2681 8407 7399
rect 3069 2640 8407 2681
rect 8807 7399 14145 7440
rect 8807 2681 13889 7399
rect 14125 2681 14145 7399
rect 8807 2640 14145 2681
rect -14145 2359 -8807 2400
rect -14145 -2359 -9063 2359
rect -8827 -2359 -8807 2359
rect -14145 -2400 -8807 -2359
rect -8407 2359 -3069 2400
rect -8407 -2359 -3325 2359
rect -3089 -2359 -3069 2359
rect -8407 -2400 -3069 -2359
rect -2669 2359 2669 2400
rect -2669 -2359 2413 2359
rect 2649 -2359 2669 2359
rect -2669 -2400 2669 -2359
rect 3069 2359 8407 2400
rect 3069 -2359 8151 2359
rect 8387 -2359 8407 2359
rect 3069 -2400 8407 -2359
rect 8807 2359 14145 2400
rect 8807 -2359 13889 2359
rect 14125 -2359 14145 2359
rect 8807 -2400 14145 -2359
rect -14145 -2681 -8807 -2640
rect -14145 -7399 -9063 -2681
rect -8827 -7399 -8807 -2681
rect -14145 -7440 -8807 -7399
rect -8407 -2681 -3069 -2640
rect -8407 -7399 -3325 -2681
rect -3089 -7399 -3069 -2681
rect -8407 -7440 -3069 -7399
rect -2669 -2681 2669 -2640
rect -2669 -7399 2413 -2681
rect 2649 -7399 2669 -2681
rect -2669 -7440 2669 -7399
rect 3069 -2681 8407 -2640
rect 3069 -7399 8151 -2681
rect 8387 -7399 8407 -2681
rect 3069 -7440 8407 -7399
rect 8807 -2681 14145 -2640
rect 8807 -7399 13889 -2681
rect 14125 -7399 14145 -2681
rect 8807 -7440 14145 -7399
rect -14145 -7721 -8807 -7680
rect -14145 -12439 -9063 -7721
rect -8827 -12439 -8807 -7721
rect -14145 -12480 -8807 -12439
rect -8407 -7721 -3069 -7680
rect -8407 -12439 -3325 -7721
rect -3089 -12439 -3069 -7721
rect -8407 -12480 -3069 -12439
rect -2669 -7721 2669 -7680
rect -2669 -12439 2413 -7721
rect 2649 -12439 2669 -7721
rect -2669 -12480 2669 -12439
rect 3069 -7721 8407 -7680
rect 3069 -12439 8151 -7721
rect 8387 -12439 8407 -7721
rect 3069 -12480 8407 -12439
rect 8807 -7721 14145 -7680
rect 8807 -12439 13889 -7721
rect 14125 -12439 14145 -7721
rect 8807 -12480 14145 -12439
<< via4 >>
rect -9063 7721 -8827 12439
rect -3325 7721 -3089 12439
rect 2413 7721 2649 12439
rect 8151 7721 8387 12439
rect 13889 7721 14125 12439
rect -9063 2681 -8827 7399
rect -3325 2681 -3089 7399
rect 2413 2681 2649 7399
rect 8151 2681 8387 7399
rect 13889 2681 14125 7399
rect -9063 -2359 -8827 2359
rect -3325 -2359 -3089 2359
rect 2413 -2359 2649 2359
rect 8151 -2359 8387 2359
rect 13889 -2359 14125 2359
rect -9063 -7399 -8827 -2681
rect -3325 -7399 -3089 -2681
rect 2413 -7399 2649 -2681
rect 8151 -7399 8387 -2681
rect 13889 -7399 14125 -2681
rect -9063 -12439 -8827 -7721
rect -3325 -12439 -3089 -7721
rect 2413 -12439 2649 -7721
rect 8151 -12439 8387 -7721
rect 13889 -12439 14125 -7721
<< mimcap2 >>
rect -14065 12360 -9425 12400
rect -14065 7800 -14025 12360
rect -9465 7800 -9425 12360
rect -14065 7760 -9425 7800
rect -8327 12360 -3687 12400
rect -8327 7800 -8287 12360
rect -3727 7800 -3687 12360
rect -8327 7760 -3687 7800
rect -2589 12360 2051 12400
rect -2589 7800 -2549 12360
rect 2011 7800 2051 12360
rect -2589 7760 2051 7800
rect 3149 12360 7789 12400
rect 3149 7800 3189 12360
rect 7749 7800 7789 12360
rect 3149 7760 7789 7800
rect 8887 12360 13527 12400
rect 8887 7800 8927 12360
rect 13487 7800 13527 12360
rect 8887 7760 13527 7800
rect -14065 7320 -9425 7360
rect -14065 2760 -14025 7320
rect -9465 2760 -9425 7320
rect -14065 2720 -9425 2760
rect -8327 7320 -3687 7360
rect -8327 2760 -8287 7320
rect -3727 2760 -3687 7320
rect -8327 2720 -3687 2760
rect -2589 7320 2051 7360
rect -2589 2760 -2549 7320
rect 2011 2760 2051 7320
rect -2589 2720 2051 2760
rect 3149 7320 7789 7360
rect 3149 2760 3189 7320
rect 7749 2760 7789 7320
rect 3149 2720 7789 2760
rect 8887 7320 13527 7360
rect 8887 2760 8927 7320
rect 13487 2760 13527 7320
rect 8887 2720 13527 2760
rect -14065 2280 -9425 2320
rect -14065 -2280 -14025 2280
rect -9465 -2280 -9425 2280
rect -14065 -2320 -9425 -2280
rect -8327 2280 -3687 2320
rect -8327 -2280 -8287 2280
rect -3727 -2280 -3687 2280
rect -8327 -2320 -3687 -2280
rect -2589 2280 2051 2320
rect -2589 -2280 -2549 2280
rect 2011 -2280 2051 2280
rect -2589 -2320 2051 -2280
rect 3149 2280 7789 2320
rect 3149 -2280 3189 2280
rect 7749 -2280 7789 2280
rect 3149 -2320 7789 -2280
rect 8887 2280 13527 2320
rect 8887 -2280 8927 2280
rect 13487 -2280 13527 2280
rect 8887 -2320 13527 -2280
rect -14065 -2760 -9425 -2720
rect -14065 -7320 -14025 -2760
rect -9465 -7320 -9425 -2760
rect -14065 -7360 -9425 -7320
rect -8327 -2760 -3687 -2720
rect -8327 -7320 -8287 -2760
rect -3727 -7320 -3687 -2760
rect -8327 -7360 -3687 -7320
rect -2589 -2760 2051 -2720
rect -2589 -7320 -2549 -2760
rect 2011 -7320 2051 -2760
rect -2589 -7360 2051 -7320
rect 3149 -2760 7789 -2720
rect 3149 -7320 3189 -2760
rect 7749 -7320 7789 -2760
rect 3149 -7360 7789 -7320
rect 8887 -2760 13527 -2720
rect 8887 -7320 8927 -2760
rect 13487 -7320 13527 -2760
rect 8887 -7360 13527 -7320
rect -14065 -7800 -9425 -7760
rect -14065 -12360 -14025 -7800
rect -9465 -12360 -9425 -7800
rect -14065 -12400 -9425 -12360
rect -8327 -7800 -3687 -7760
rect -8327 -12360 -8287 -7800
rect -3727 -12360 -3687 -7800
rect -8327 -12400 -3687 -12360
rect -2589 -7800 2051 -7760
rect -2589 -12360 -2549 -7800
rect 2011 -12360 2051 -7800
rect -2589 -12400 2051 -12360
rect 3149 -7800 7789 -7760
rect 3149 -12360 3189 -7800
rect 7749 -12360 7789 -7800
rect 3149 -12400 7789 -12360
rect 8887 -7800 13527 -7760
rect 8887 -12360 8927 -7800
rect 13487 -12360 13527 -7800
rect 8887 -12400 13527 -12360
<< mimcap2contact >>
rect -14025 7800 -9465 12360
rect -8287 7800 -3727 12360
rect -2549 7800 2011 12360
rect 3189 7800 7749 12360
rect 8927 7800 13487 12360
rect -14025 2760 -9465 7320
rect -8287 2760 -3727 7320
rect -2549 2760 2011 7320
rect 3189 2760 7749 7320
rect 8927 2760 13487 7320
rect -14025 -2280 -9465 2280
rect -8287 -2280 -3727 2280
rect -2549 -2280 2011 2280
rect 3189 -2280 7749 2280
rect 8927 -2280 13487 2280
rect -14025 -7320 -9465 -2760
rect -8287 -7320 -3727 -2760
rect -2549 -7320 2011 -2760
rect 3189 -7320 7749 -2760
rect 8927 -7320 13487 -2760
rect -14025 -12360 -9465 -7800
rect -8287 -12360 -3727 -7800
rect -2549 -12360 2011 -7800
rect 3189 -12360 7749 -7800
rect 8927 -12360 13487 -7800
<< metal5 >>
rect -11905 12384 -11585 12600
rect -9105 12439 -8785 12600
rect -14049 12360 -9441 12384
rect -14049 7800 -14025 12360
rect -9465 7800 -9441 12360
rect -14049 7776 -9441 7800
rect -11905 7344 -11585 7776
rect -9105 7721 -9063 12439
rect -8827 7721 -8785 12439
rect -6167 12384 -5847 12600
rect -3367 12439 -3047 12600
rect -8311 12360 -3703 12384
rect -8311 7800 -8287 12360
rect -3727 7800 -3703 12360
rect -8311 7776 -3703 7800
rect -9105 7399 -8785 7721
rect -14049 7320 -9441 7344
rect -14049 2760 -14025 7320
rect -9465 2760 -9441 7320
rect -14049 2736 -9441 2760
rect -11905 2304 -11585 2736
rect -9105 2681 -9063 7399
rect -8827 2681 -8785 7399
rect -6167 7344 -5847 7776
rect -3367 7721 -3325 12439
rect -3089 7721 -3047 12439
rect -429 12384 -109 12600
rect 2371 12439 2691 12600
rect -2573 12360 2035 12384
rect -2573 7800 -2549 12360
rect 2011 7800 2035 12360
rect -2573 7776 2035 7800
rect -3367 7399 -3047 7721
rect -8311 7320 -3703 7344
rect -8311 2760 -8287 7320
rect -3727 2760 -3703 7320
rect -8311 2736 -3703 2760
rect -9105 2359 -8785 2681
rect -14049 2280 -9441 2304
rect -14049 -2280 -14025 2280
rect -9465 -2280 -9441 2280
rect -14049 -2304 -9441 -2280
rect -11905 -2736 -11585 -2304
rect -9105 -2359 -9063 2359
rect -8827 -2359 -8785 2359
rect -6167 2304 -5847 2736
rect -3367 2681 -3325 7399
rect -3089 2681 -3047 7399
rect -429 7344 -109 7776
rect 2371 7721 2413 12439
rect 2649 7721 2691 12439
rect 5309 12384 5629 12600
rect 8109 12439 8429 12600
rect 3165 12360 7773 12384
rect 3165 7800 3189 12360
rect 7749 7800 7773 12360
rect 3165 7776 7773 7800
rect 2371 7399 2691 7721
rect -2573 7320 2035 7344
rect -2573 2760 -2549 7320
rect 2011 2760 2035 7320
rect -2573 2736 2035 2760
rect -3367 2359 -3047 2681
rect -8311 2280 -3703 2304
rect -8311 -2280 -8287 2280
rect -3727 -2280 -3703 2280
rect -8311 -2304 -3703 -2280
rect -9105 -2681 -8785 -2359
rect -14049 -2760 -9441 -2736
rect -14049 -7320 -14025 -2760
rect -9465 -7320 -9441 -2760
rect -14049 -7344 -9441 -7320
rect -11905 -7776 -11585 -7344
rect -9105 -7399 -9063 -2681
rect -8827 -7399 -8785 -2681
rect -6167 -2736 -5847 -2304
rect -3367 -2359 -3325 2359
rect -3089 -2359 -3047 2359
rect -429 2304 -109 2736
rect 2371 2681 2413 7399
rect 2649 2681 2691 7399
rect 5309 7344 5629 7776
rect 8109 7721 8151 12439
rect 8387 7721 8429 12439
rect 11047 12384 11367 12600
rect 13847 12439 14167 12600
rect 8903 12360 13511 12384
rect 8903 7800 8927 12360
rect 13487 7800 13511 12360
rect 8903 7776 13511 7800
rect 8109 7399 8429 7721
rect 3165 7320 7773 7344
rect 3165 2760 3189 7320
rect 7749 2760 7773 7320
rect 3165 2736 7773 2760
rect 2371 2359 2691 2681
rect -2573 2280 2035 2304
rect -2573 -2280 -2549 2280
rect 2011 -2280 2035 2280
rect -2573 -2304 2035 -2280
rect -3367 -2681 -3047 -2359
rect -8311 -2760 -3703 -2736
rect -8311 -7320 -8287 -2760
rect -3727 -7320 -3703 -2760
rect -8311 -7344 -3703 -7320
rect -9105 -7721 -8785 -7399
rect -14049 -7800 -9441 -7776
rect -14049 -12360 -14025 -7800
rect -9465 -12360 -9441 -7800
rect -14049 -12384 -9441 -12360
rect -11905 -12600 -11585 -12384
rect -9105 -12439 -9063 -7721
rect -8827 -12439 -8785 -7721
rect -6167 -7776 -5847 -7344
rect -3367 -7399 -3325 -2681
rect -3089 -7399 -3047 -2681
rect -429 -2736 -109 -2304
rect 2371 -2359 2413 2359
rect 2649 -2359 2691 2359
rect 5309 2304 5629 2736
rect 8109 2681 8151 7399
rect 8387 2681 8429 7399
rect 11047 7344 11367 7776
rect 13847 7721 13889 12439
rect 14125 7721 14167 12439
rect 13847 7399 14167 7721
rect 8903 7320 13511 7344
rect 8903 2760 8927 7320
rect 13487 2760 13511 7320
rect 8903 2736 13511 2760
rect 8109 2359 8429 2681
rect 3165 2280 7773 2304
rect 3165 -2280 3189 2280
rect 7749 -2280 7773 2280
rect 3165 -2304 7773 -2280
rect 2371 -2681 2691 -2359
rect -2573 -2760 2035 -2736
rect -2573 -7320 -2549 -2760
rect 2011 -7320 2035 -2760
rect -2573 -7344 2035 -7320
rect -3367 -7721 -3047 -7399
rect -8311 -7800 -3703 -7776
rect -8311 -12360 -8287 -7800
rect -3727 -12360 -3703 -7800
rect -8311 -12384 -3703 -12360
rect -9105 -12600 -8785 -12439
rect -6167 -12600 -5847 -12384
rect -3367 -12439 -3325 -7721
rect -3089 -12439 -3047 -7721
rect -429 -7776 -109 -7344
rect 2371 -7399 2413 -2681
rect 2649 -7399 2691 -2681
rect 5309 -2736 5629 -2304
rect 8109 -2359 8151 2359
rect 8387 -2359 8429 2359
rect 11047 2304 11367 2736
rect 13847 2681 13889 7399
rect 14125 2681 14167 7399
rect 13847 2359 14167 2681
rect 8903 2280 13511 2304
rect 8903 -2280 8927 2280
rect 13487 -2280 13511 2280
rect 8903 -2304 13511 -2280
rect 8109 -2681 8429 -2359
rect 3165 -2760 7773 -2736
rect 3165 -7320 3189 -2760
rect 7749 -7320 7773 -2760
rect 3165 -7344 7773 -7320
rect 2371 -7721 2691 -7399
rect -2573 -7800 2035 -7776
rect -2573 -12360 -2549 -7800
rect 2011 -12360 2035 -7800
rect -2573 -12384 2035 -12360
rect -3367 -12600 -3047 -12439
rect -429 -12600 -109 -12384
rect 2371 -12439 2413 -7721
rect 2649 -12439 2691 -7721
rect 5309 -7776 5629 -7344
rect 8109 -7399 8151 -2681
rect 8387 -7399 8429 -2681
rect 11047 -2736 11367 -2304
rect 13847 -2359 13889 2359
rect 14125 -2359 14167 2359
rect 13847 -2681 14167 -2359
rect 8903 -2760 13511 -2736
rect 8903 -7320 8927 -2760
rect 13487 -7320 13511 -2760
rect 8903 -7344 13511 -7320
rect 8109 -7721 8429 -7399
rect 3165 -7800 7773 -7776
rect 3165 -12360 3189 -7800
rect 7749 -12360 7773 -7800
rect 3165 -12384 7773 -12360
rect 2371 -12600 2691 -12439
rect 5309 -12600 5629 -12384
rect 8109 -12439 8151 -7721
rect 8387 -12439 8429 -7721
rect 11047 -7776 11367 -7344
rect 13847 -7399 13889 -2681
rect 14125 -7399 14167 -2681
rect 13847 -7721 14167 -7399
rect 8903 -7800 13511 -7776
rect 8903 -12360 8927 -7800
rect 13487 -12360 13511 -7800
rect 8903 -12384 13511 -12360
rect 8109 -12600 8429 -12439
rect 11047 -12600 11367 -12384
rect 13847 -12439 13889 -7721
rect 14125 -12439 14167 -7721
rect 13847 -12600 14167 -12439
<< properties >>
string FIXED_BBOX 8807 7680 13607 12480
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.2 l 23.2 val 1.094k carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
