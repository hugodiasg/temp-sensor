magic
tech sky130A
timestamp 1644594744
<< pwell >>
rect -139 -564 139 564
<< mvnmos >>
rect -25 -435 25 435
<< mvndiff >>
rect -54 429 -25 435
rect -54 -429 -48 429
rect -31 -429 -25 429
rect -54 -435 -25 -429
rect 25 429 54 435
rect 25 -429 31 429
rect 48 -429 54 429
rect 25 -435 54 -429
<< mvndiffc >>
rect -48 -429 -31 429
rect 31 -429 48 429
<< mvpsubdiff >>
rect -121 540 121 546
rect -121 523 -67 540
rect 67 523 121 540
rect -121 517 121 523
rect -121 492 -92 517
rect -121 -492 -115 492
rect -98 -492 -92 492
rect 92 492 121 517
rect -121 -517 -92 -492
rect 92 -492 98 492
rect 115 -492 121 492
rect 92 -517 121 -492
rect -121 -523 121 -517
rect -121 -540 -67 -523
rect 67 -540 121 -523
rect -121 -546 121 -540
<< mvpsubdiffcont >>
rect -67 523 67 540
rect -115 -492 -98 492
rect 98 -492 115 492
rect -67 -540 67 -523
<< poly >>
rect -25 471 25 479
rect -25 454 -17 471
rect 17 454 25 471
rect -25 435 25 454
rect -25 -454 25 -435
rect -25 -471 -17 -454
rect 17 -471 25 -454
rect -25 -479 25 -471
<< polycont >>
rect -17 454 17 471
rect -17 -471 17 -454
<< locali >>
rect -115 492 -98 540
rect 98 492 115 540
rect -25 454 -17 471
rect 17 454 25 471
rect -48 429 -31 437
rect -48 -437 -31 -429
rect 31 429 48 437
rect 31 -437 48 -429
rect -25 -471 -17 -454
rect 17 -471 25 -454
rect -115 -523 -98 -492
rect 98 -523 115 -492
rect -115 -540 -67 -523
rect 67 -540 115 -523
<< viali >>
rect -98 523 -67 540
rect -67 523 67 540
rect 67 523 98 540
rect -17 454 17 471
rect -48 -429 -31 429
rect 31 -429 48 429
rect -17 -471 17 -454
<< metal1 >>
rect -104 540 104 543
rect -104 523 -98 540
rect 98 523 104 540
rect -104 520 104 523
rect -23 471 23 474
rect -23 454 -17 471
rect 17 454 23 471
rect -23 451 23 454
rect -51 429 -28 435
rect -51 -429 -48 429
rect -31 -429 -28 429
rect -51 -435 -28 -429
rect 28 429 51 435
rect 28 -429 31 429
rect 48 -429 51 429
rect 28 -435 51 -429
rect -23 -454 23 -451
rect -23 -471 -17 -454
rect 17 -471 23 -454
rect -23 -474 23 -471
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -106 -531 106 531
string parameters w 8.7 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
string library sky130
<< end >>
