magic
tech sky130A
magscale 1 2
timestamp 1646019513
<< metal4 >>
rect -2611 7655 2611 7696
rect -2611 2673 2355 7655
rect 2591 2673 2611 7655
rect -2611 2632 2611 2673
rect -2611 2491 2611 2532
rect -2611 -2491 2355 2491
rect 2591 -2491 2611 2491
rect -2611 -2532 2611 -2491
rect -2611 -2673 2611 -2632
rect -2611 -7655 2355 -2673
rect 2591 -7655 2611 -2673
rect -2611 -7696 2611 -7655
<< via4 >>
rect 2355 2673 2591 7655
rect 2355 -2491 2591 2491
rect 2355 -7655 2591 -2673
<< mimcap2 >>
rect -2511 7556 2353 7596
rect -2511 2772 -1993 7556
rect 1835 2772 2353 7556
rect -2511 2732 2353 2772
rect -2511 2392 2353 2432
rect -2511 -2392 -1993 2392
rect 1835 -2392 2353 2392
rect -2511 -2432 2353 -2392
rect -2511 -2772 2353 -2732
rect -2511 -7556 -1993 -2772
rect 1835 -7556 2353 -2772
rect -2511 -7596 2353 -7556
<< mimcap2contact >>
rect -1993 2772 1835 7556
rect -1993 -2392 1835 2392
rect -1993 -7556 1835 -2772
<< metal5 >>
rect -239 7580 81 7746
rect 2313 7655 2633 7746
rect -2017 7556 1859 7580
rect -2017 2772 -1993 7556
rect 1835 2772 1859 7556
rect -2017 2748 1859 2772
rect -239 2416 81 2748
rect 2313 2673 2355 7655
rect 2591 2673 2633 7655
rect 2313 2491 2633 2673
rect -2017 2392 1859 2416
rect -2017 -2392 -1993 2392
rect 1835 -2392 1859 2392
rect -2017 -2416 1859 -2392
rect -239 -2748 81 -2416
rect 2313 -2491 2355 2491
rect 2591 -2491 2633 2491
rect 2313 -2673 2633 -2491
rect -2017 -2772 1859 -2748
rect -2017 -7556 -1993 -2772
rect 1835 -7556 1859 -2772
rect -2017 -7580 1859 -7556
rect -239 -7746 81 -7580
rect 2313 -7655 2355 -2673
rect 2591 -7655 2633 -2673
rect 2313 -7746 2633 -7655
<< properties >>
string FIXED_BBOX -2611 2632 2453 7696
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.315 l 24.315 val 1.2k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
