magic
tech sky130A
magscale 1 2
timestamp 1644161670
<< error_p >>
rect 1919 2716 2003 7484
rect 1919 -2384 2003 2384
rect 1919 -7484 2003 -2716
rect 2239 -7650 2323 7650
rect 2559 2599 2643 2821
rect 2559 2279 2643 2501
rect 2559 -2501 2643 -2279
rect 2559 -2821 2643 -2599
<< metal4 >>
rect -2621 7559 2621 7600
rect -2621 2641 2365 7559
rect 2601 2641 2621 7559
rect -2621 2600 2621 2641
rect -2621 2459 2621 2500
rect -2621 -2459 2365 2459
rect 2601 -2459 2621 2459
rect -2621 -2500 2621 -2459
rect -2621 -2641 2621 -2600
rect -2621 -7559 2365 -2641
rect 2601 -7559 2621 -2641
rect -2621 -7600 2621 -7559
<< via4 >>
rect 2365 2641 2601 7559
rect 2365 -2459 2601 2459
rect 2365 -7559 2601 -2641
<< mimcap2 >>
rect -2521 7460 2279 7500
rect -2521 2740 -2221 7460
rect 1979 2740 2279 7460
rect -2521 2700 2279 2740
rect -2521 2360 2279 2400
rect -2521 -2360 -2221 2360
rect 1979 -2360 2279 2360
rect -2521 -2400 2279 -2360
rect -2521 -2740 2279 -2700
rect -2521 -7460 -2221 -2740
rect 1979 -7460 2279 -2740
rect -2521 -7500 2279 -7460
<< mimcap2contact >>
rect -2221 2740 1979 7460
rect -2221 -2360 1979 2360
rect -2221 -7460 1979 -2740
<< metal5 >>
rect -281 7484 39 7650
rect 2239 7601 2559 7650
rect 2239 7559 2643 7601
rect -2245 7460 2003 7484
rect -2245 2740 -2221 7460
rect 1979 2740 2003 7460
rect -2245 2716 2003 2740
rect -281 2384 39 2716
rect 2239 2641 2365 7559
rect 2601 2641 2643 7559
rect 2239 2599 2643 2641
rect 2239 2501 2559 2599
rect 2239 2459 2643 2501
rect -2245 2360 2003 2384
rect -2245 -2360 -2221 2360
rect 1979 -2360 2003 2360
rect -2245 -2384 2003 -2360
rect -281 -2716 39 -2384
rect 2239 -2459 2365 2459
rect 2601 -2459 2643 2459
rect 2239 -2501 2643 -2459
rect 2239 -2599 2559 -2501
rect 2239 -2641 2643 -2599
rect -2245 -2740 2003 -2716
rect -2245 -7460 -2221 -2740
rect 1979 -7460 2003 -2740
rect -2245 -7484 2003 -7460
rect -281 -7650 39 -7484
rect 2239 -7559 2365 -2641
rect 2601 -7559 2643 -2641
rect 2239 -7601 2643 -7559
rect 2239 -7650 2559 -7601
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2621 2600 2379 7600
string parameters w 24.0 l 24.0 val 1.17k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 89
string library sky130
<< end >>
