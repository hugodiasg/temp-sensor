magic
tech sky130A
magscale 1 2
timestamp 1645034691
<< metal4 >>
rect -2639 7739 2639 7780
rect -2639 2701 2383 7739
rect 2619 2701 2639 7739
rect -2639 2660 2639 2701
rect -2639 2519 2639 2560
rect -2639 -2519 2383 2519
rect 2619 -2519 2639 2519
rect -2639 -2560 2639 -2519
rect -2639 -2701 2639 -2660
rect -2639 -7739 2383 -2701
rect 2619 -7739 2639 -2701
rect -2639 -7780 2639 -7739
<< via4 >>
rect 2383 2701 2619 7739
rect 2383 -2519 2619 2519
rect 2383 -7739 2619 -2701
<< mimcap2 >>
rect -2539 7640 2381 7680
rect -2539 2800 -2015 7640
rect 1857 2800 2381 7640
rect -2539 2760 2381 2800
rect -2539 2420 2381 2460
rect -2539 -2420 -2015 2420
rect 1857 -2420 2381 2420
rect -2539 -2460 2381 -2420
rect -2539 -2800 2381 -2760
rect -2539 -7640 -2015 -2800
rect 1857 -7640 2381 -2800
rect -2539 -7680 2381 -7640
<< mimcap2contact >>
rect -2015 2800 1857 7640
rect -2015 -2420 1857 2420
rect -2015 -7640 1857 -2800
<< metal5 >>
rect -239 7664 81 7830
rect 2341 7739 2661 7830
rect -2039 7640 1881 7664
rect -2039 2800 -2015 7640
rect 1857 2800 1881 7640
rect -2039 2776 1881 2800
rect -239 2444 81 2776
rect 2341 2701 2383 7739
rect 2619 2701 2661 7739
rect 2341 2519 2661 2701
rect -2039 2420 1881 2444
rect -2039 -2420 -2015 2420
rect 1857 -2420 1881 2420
rect -2039 -2444 1881 -2420
rect -239 -2776 81 -2444
rect 2341 -2519 2383 2519
rect 2619 -2519 2661 2519
rect 2341 -2701 2661 -2519
rect -2039 -2800 1881 -2776
rect -2039 -7640 -2015 -2800
rect 1857 -7640 1881 -2800
rect -2039 -7664 1881 -7640
rect -239 -7830 81 -7664
rect 2341 -7739 2383 -2701
rect 2619 -7739 2661 -2701
rect 2341 -7830 2661 -7739
<< properties >>
string FIXED_BBOX -2639 2660 2481 7780
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.6 l 24.6 val 1.229k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
