magic
tech sky130A
magscale 1 2
timestamp 1645495691
<< metal4 >>
rect -3080 12113 3080 12154
rect -3080 6193 2824 12113
rect 3060 6193 3080 12113
rect -3080 6152 3080 6193
rect -3080 6011 3080 6052
rect -3080 91 2824 6011
rect 3060 91 3080 6011
rect -3080 50 3080 91
rect -3080 -91 3080 -50
rect -3080 -6011 2824 -91
rect 3060 -6011 3080 -91
rect -3080 -6052 3080 -6011
rect -3080 -6193 3080 -6152
rect -3080 -12113 2824 -6193
rect 3060 -12113 3080 -6193
rect -3080 -12154 3080 -12113
<< via4 >>
rect 2824 6193 3060 12113
rect 2824 91 3060 6011
rect 2824 -6011 3060 -91
rect 2824 -12113 3060 -6193
<< mimcap2 >>
rect -2980 12014 2822 12054
rect -2980 6292 -2368 12014
rect 2210 6292 2822 12014
rect -2980 6252 2822 6292
rect -2980 5912 2822 5952
rect -2980 190 -2368 5912
rect 2210 190 2822 5912
rect -2980 150 2822 190
rect -2980 -190 2822 -150
rect -2980 -5912 -2368 -190
rect 2210 -5912 2822 -190
rect -2980 -5952 2822 -5912
rect -2980 -6292 2822 -6252
rect -2980 -12014 -2368 -6292
rect 2210 -12014 2822 -6292
rect -2980 -12054 2822 -12014
<< mimcap2contact >>
rect -2368 6292 2210 12014
rect -2368 190 2210 5912
rect -2368 -5912 2210 -190
rect -2368 -12014 2210 -6292
<< metal5 >>
rect -239 12038 81 12204
rect 2782 12113 3102 12204
rect -2392 12014 2234 12038
rect -2392 6292 -2368 12014
rect 2210 6292 2234 12014
rect -2392 6268 2234 6292
rect -239 5936 81 6268
rect 2782 6193 2824 12113
rect 3060 6193 3102 12113
rect 2782 6011 3102 6193
rect -2392 5912 2234 5936
rect -2392 190 -2368 5912
rect 2210 190 2234 5912
rect -2392 166 2234 190
rect -239 -166 81 166
rect 2782 91 2824 6011
rect 3060 91 3102 6011
rect 2782 -91 3102 91
rect -2392 -190 2234 -166
rect -2392 -5912 -2368 -190
rect 2210 -5912 2234 -190
rect -2392 -5936 2234 -5912
rect -239 -6268 81 -5936
rect 2782 -6011 2824 -91
rect 3060 -6011 3102 -91
rect 2782 -6193 3102 -6011
rect -2392 -6292 2234 -6268
rect -2392 -12014 -2368 -6292
rect 2210 -12014 2234 -6292
rect -2392 -12038 2234 -12014
rect -239 -12204 81 -12038
rect 2782 -12113 2824 -6193
rect 3060 -12113 3102 -6193
rect 2782 -12204 3102 -12113
<< properties >>
string FIXED_BBOX -3080 6152 2922 12154
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 29.008 l 29.008 val 1.704k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
