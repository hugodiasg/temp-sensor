* NGSPICE file created from ask-modulator.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN w_n201_n1098# a_n35_500# a_n35_n932#
X0 a_n35_n932# a_n35_500# w_n201_n1098# sky130_fd_pr__res_xhigh_po_0p35 l=5e+06u
C0 a_n35_n932# w_n201_n1098# 1.08fF
C1 a_n35_500# w_n201_n1098# 1.08fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_9XH3MC c2_n2414_n7305# m4_n2514_n7405# VSUBS
X0 c2_n2414_n7305# m4_n2514_n7405# sky130_fd_pr__cap_mim_m3_2 l=2.335e+07u w=2.335e+07u
X1 c2_n2414_n7305# m4_n2514_n7405# sky130_fd_pr__cap_mim_m3_2 l=2.335e+07u w=2.335e+07u
X2 c2_n2414_n7305# m4_n2514_n7405# sky130_fd_pr__cap_mim_m3_2 l=2.335e+07u w=2.335e+07u
C0 m4_n2514_n7405# c2_n2414_n7305# 109.41fF
C1 c2_n2414_n7305# VSUBS 0.26fF
C2 m4_n2514_n7405# VSUBS 28.83fF
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PWYS4E a_n108_n870# a_n50_n958# w_n278_n1128#
+ a_50_n870#
X0 a_50_n870# a_n50_n958# a_n108_n870# w_n278_n1128# sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=8.7e+06u l=500000u
C0 a_50_n870# a_n108_n870# 1.03fF
C1 a_50_n870# w_n278_n1128# 0.84fF
C2 a_n108_n870# w_n278_n1128# 0.84fF
C3 a_n50_n958# w_n278_n1128# 0.52fF
.ends

.subckt ask-modulator in out vd gnd
Xsky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0 gnd vd out sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN
Xsky130_fd_pr__cap_mim_m3_2_9XH3MC_0 vd out gnd sky130_fd_pr__cap_mim_m3_2_9XH3MC
Xsky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5_PWYS4E
X0 vd.t1 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
X1 vd.t2 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
X2 vd.t0 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 out vd sky130_fd_pr__res_generic_m4 w=6e+06u l=900000u
X3 gnd in.t0 out gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=0u l=0u
R1 vd vd.t1 2.666
R2 vd.t0 vd.t2 0.066
R3 vd.t1 vd.t0 0.066
R4 in in.t0 448.598
C0 out in 0.46fF
C1 out vd 0.14fF
C2 m4_11480_14620# gnd 0.11fF $ **FLOATING
C3 in.t0 gnd 0.45fF
C4 vd.t2 gnd 25.05fF
C5 vd.t0 gnd 25.12fF
C6 vd.t1 gnd 173.47fF
C7 out gnd 200.74fF
C8 in gnd 5.53fF
C9 vd gnd 136.30fF
.ends

