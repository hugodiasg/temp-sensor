magic
tech sky130A
magscale 1 2
timestamp 1646008289
<< mvpsubdiff >>
rect 406200 555400 408200 555424
rect 406200 552976 408200 553000
<< mvpsubdiffcont >>
rect 406200 553000 408200 555400
<< locali >>
rect 406200 555400 408200 555416
rect 406200 552984 408200 553000
<< viali >>
rect 406200 553000 408200 555400
<< metal1 >>
rect 414500 591600 430000 592000
rect 414500 587000 415200 591600
rect 404800 581600 415200 587000
rect 414500 577200 415200 581600
rect 429600 577200 430000 591600
rect 414500 576600 430000 577200
rect 404800 557800 413600 558000
rect 404800 555800 410400 557800
rect 413400 555800 413600 557800
rect 404800 555600 413600 555800
rect 406000 555400 408400 555600
rect 406000 553000 406200 555400
rect 408200 553000 408400 555400
rect 406000 552800 408400 553000
rect 410400 530400 430600 531000
rect 410400 526400 411000 530400
rect 404800 521000 411000 526400
rect 410400 515600 411000 521000
rect 430200 515600 430600 530400
rect 410400 515400 430600 515600
<< via1 >>
rect 415200 577200 429600 591600
rect 410400 555800 413400 557800
rect 411000 515600 430200 530400
<< metal2 >>
rect 414500 591600 430000 592000
rect 414500 577200 415200 591600
rect 429600 577200 430000 591600
rect 414500 576600 430000 577200
rect 408000 557800 413600 558000
rect 408000 555800 410400 557800
rect 413400 555800 413600 557800
rect 408000 555600 413600 555800
rect 410400 530400 430600 531000
rect 410400 515600 411000 530400
rect 430200 515600 430600 530400
rect 410400 515400 430600 515600
<< via2 >>
rect 415200 577200 429600 591600
rect 410400 555800 413400 557800
rect 411000 515600 430200 530400
<< metal3 >>
rect 414500 591600 430000 592000
rect 414500 577200 415200 591600
rect 429600 577200 430000 591600
rect 414500 576600 430000 577200
rect 408000 557800 413600 558000
rect 408000 555800 410400 557800
rect 413400 555800 413600 557800
rect 408000 555600 413600 555800
rect 410400 530400 430600 531000
rect 410400 515600 411000 530400
rect 430200 515600 430600 530400
rect 410400 515400 430600 515600
<< via3 >>
rect 415200 577200 429600 591600
rect 410400 555800 413400 557800
rect 411000 515600 430200 530400
<< metal4 >>
rect 414500 591600 430000 592000
rect 414500 577200 415200 591600
rect 429600 577200 430000 591600
rect 414500 576600 430000 577200
rect 415600 558000 418600 562200
rect 421200 558000 424200 562200
rect 426600 558000 429600 562200
rect 408000 557800 429600 558000
rect 408000 555800 410400 557800
rect 413400 555800 429600 557800
rect 408000 555600 429600 555800
rect 410200 552600 413200 555600
rect 415600 552000 418600 555600
rect 421200 551800 424200 555600
rect 426600 552400 429600 555600
rect 410400 530400 430600 531000
rect 410400 515600 411000 530400
rect 430200 515600 430600 530400
rect 410400 515400 430600 515600
<< via4 >>
rect 415200 577200 429600 591600
rect 411000 515600 430200 530400
<< metal5 >>
rect 414500 591600 430600 592000
rect 414500 577200 415200 591600
rect 429600 577200 430600 591600
rect 414500 576600 430600 577200
rect 432000 576600 447400 592000
rect 415000 570400 418000 576600
rect 421000 570400 424000 576600
rect 425800 570600 428800 576600
rect 410400 531000 412800 536000
rect 415600 531000 418600 536000
rect 421400 531000 424400 536000
rect 427000 531000 430000 536400
rect 410400 530400 430400 531000
rect 410400 515600 411000 530400
rect 430200 515600 430400 530400
rect 410400 515400 430400 515600
<< rm5 >>
rect 430600 576600 432000 592000
use l0  l0_0
timestamp 1645758648
transform 1 0 0 0 1 0
box 418100 432000 592000 592000
use sky130_fd_pr__cap_mim_m3_2_3YFQRG  sky130_fd_pr__cap_mim_m3_2_3YFQRG_0
timestamp 1645800166
transform 1 0 411354 0 1 544267
box -2675 -10584 2697 10584
use sky130_fd_pr__cap_mim_m3_2_3YFQRG  sky130_fd_pr__cap_mim_m3_2_3YFQRG_1
timestamp 1645800166
transform 1 0 417289 0 1 544461
box -2675 -10584 2697 10584
use sky130_fd_pr__cap_mim_m3_2_3YFQRG  sky130_fd_pr__cap_mim_m3_2_3YFQRG_2
timestamp 1645800166
transform 1 0 423089 0 1 544411
box -2675 -10584 2697 10584
use sky130_fd_pr__cap_mim_m3_2_3YFQRG  sky130_fd_pr__cap_mim_m3_2_3YFQRG_3
timestamp 1645800166
transform 1 0 428732 0 1 544329
box -2675 -10584 2697 10584
use sky130_fd_pr__cap_mim_m3_2_93FFAE  sky130_fd_pr__cap_mim_m3_2_93FFAE_0
timestamp 1645800166
transform 1 0 417022 0 1 566779
box -2622 -7779 2644 7779
use sky130_fd_pr__cap_mim_m3_2_93FFAE  sky130_fd_pr__cap_mim_m3_2_93FFAE_1
timestamp 1645800166
transform 1 0 422544 0 1 566801
box -2622 -7779 2644 7779
use sky130_fd_pr__cap_mim_m3_2_93FFAE  sky130_fd_pr__cap_mim_m3_2_93FFAE_2
timestamp 1645800166
transform 1 0 428022 0 1 566779
box -2622 -7779 2644 7779
<< labels >>
flabel metal1 405400 555800 407200 557600 0 FreeSans 1600 0 0 0 gnd
port 2 nsew
flabel metal1 406000 583600 407800 585400 0 FreeSans 1600 0 0 0 in
port 5 nsew
flabel metal1 405600 522400 408000 525000 0 FreeSans 1600 0 0 0 out
port 4 nsew
<< end >>
