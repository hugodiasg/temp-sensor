** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer.sch
.subckt impedance-transformer gnd in out
*.PININFO gnd:B in:B out:B
XC0 in gnd sky130_fd_pr__cap_mim_m3_2 W=21.5 L=21.5 MF=9 m=9
XC1 out gnd sky130_fd_pr__cap_mim_m3_2 W=26.643 L=26.643 MF=12 m=12
.ends
.end
