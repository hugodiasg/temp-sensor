magic
tech sky130A
magscale 1 2
timestamp 1661710099
<< metal1 >>
rect 3512 9225 3688 9488
rect 3512 9095 8460 9225
rect 3512 9072 3688 9095
rect -410 7800 200 7820
rect -410 7630 10 7800
rect 190 7630 200 7800
rect 8330 7720 8460 9095
rect -410 7620 200 7630
rect -400 6720 200 6920
rect 6700 6720 8480 6920
rect 8280 5990 8470 6000
rect 8280 5810 8290 5990
rect 8460 5810 8470 5990
rect 16465 5840 16865 5950
rect 8280 5800 8470 5810
rect -380 5480 200 5680
rect 10170 5060 10180 5200
rect 10320 5060 10330 5200
rect -380 4810 230 4820
rect -380 4630 -10 4810
rect 220 4630 230 4810
rect -380 4620 230 4630
<< via1 >>
rect 10 7630 190 7800
rect 8290 5810 8460 5990
rect 10180 5060 10320 5200
rect -10 4630 220 4810
<< metal2 >>
rect -10 7800 200 7820
rect -10 7630 10 7800
rect 190 7630 200 7800
rect -10 7620 200 7630
rect 8280 5990 8470 6000
rect 8280 5810 8290 5990
rect 8460 5810 8470 5990
rect 8280 5800 8470 5810
rect 10170 5200 10340 5210
rect 10170 5060 10180 5200
rect 10320 5060 10340 5200
rect 10170 5050 10340 5060
rect -20 4810 230 4820
rect -20 4630 -10 4810
rect 220 4630 230 4810
rect -20 4620 230 4630
<< via2 >>
rect 10 7630 190 7800
rect 8290 5810 8460 5990
rect 10180 5060 10320 5200
rect -10 4630 220 4810
<< metal3 >>
rect -10 7800 7645 7830
rect -10 7630 10 7800
rect 190 7630 7645 7800
rect -10 7620 7645 7630
rect 1005 6145 6035 6315
rect -20 4810 230 4820
rect -20 4630 -10 4810
rect 220 4795 230 4810
rect 1005 4795 1175 6145
rect 5865 5220 6035 6145
rect 7435 6005 7645 7620
rect 7435 5990 8475 6005
rect 7435 5810 8290 5990
rect 8460 5810 8475 5990
rect 7435 5795 8475 5810
rect 5865 5200 10330 5220
rect 5865 5060 10180 5200
rect 10320 5060 10330 5200
rect 5865 5050 10330 5060
rect 220 4630 1175 4795
rect -20 4625 1175 4630
rect -20 4620 230 4625
use buffer  buffer_0 ~/projects-sky130/temp-sensor/amp-op/mag/buffer/mag
timestamp 1661709424
transform 1 0 -5545 0 1 3610
box 13875 1430 22120 4948
use ota  ota_0 ~/projects-sky130/temp-sensor/amp-op/mag/ota
timestamp 1657059275
transform 1 0 1040 0 1 -3600
box -1040 3600 6114 12960
<< labels >>
flabel metal1 3520 9350 3680 9480 0 FreeSans 3200 0 0 0 vd
port 0 nsew
flabel metal1 -390 7640 -230 7770 0 FreeSans 3200 0 0 0 ib
port 1 nsew
flabel metal1 -390 6740 -230 6870 0 FreeSans 3200 0 0 0 in2
port 2 nsew
flabel metal1 -370 5500 -210 5630 0 FreeSans 3200 0 0 0 in1
port 3 nsew
flabel metal1 -350 4640 -190 4770 0 FreeSans 3200 0 0 0 vs
port 4 nsew
flabel metal1 16740 5850 16850 5940 0 FreeSans 3200 0 0 0 out
port 5 nsew
<< end >>
