magic
tech sky130A
magscale 1 2
timestamp 1700177945
<< nwell >>
rect 9767 2960 16933 3433
rect 9767 2940 14840 2960
rect 14900 2940 16933 2960
rect 9767 2747 16933 2940
<< pwell >>
rect 9820 1860 16212 2480
rect 9900 1020 16680 1640
<< psubdiff >>
rect 9856 2410 9952 2444
rect 16080 2410 16176 2444
rect 9856 2348 9890 2410
rect 9856 1930 9890 1992
rect 16142 2348 16176 2410
rect 16142 1930 16176 1992
rect 9856 1896 9952 1930
rect 16080 1896 16176 1930
rect 9936 1570 10032 1604
rect 16560 1570 16656 1604
rect 9936 1508 9970 1570
rect 9936 1090 9970 1152
rect 16622 1508 16656 1570
rect 16622 1090 16656 1152
rect 9936 1056 10032 1090
rect 16560 1056 16656 1090
<< nsubdiff >>
rect 9803 3363 9863 3397
rect 16837 3363 16897 3397
rect 9803 3337 9837 3363
rect 9803 2817 9837 2843
rect 16863 3337 16897 3363
rect 16863 2817 16897 2843
rect 9803 2783 9863 2817
rect 16837 2783 16897 2817
<< psubdiffcont >>
rect 9952 2410 16080 2444
rect 9856 1992 9890 2348
rect 16142 1992 16176 2348
rect 9952 1896 16080 1930
rect 10032 1570 16560 1604
rect 9936 1152 9970 1508
rect 16622 1152 16656 1508
rect 10032 1056 16560 1090
<< nsubdiffcont >>
rect 9863 3363 16837 3397
rect 9803 2843 9837 3337
rect 16863 2843 16897 3337
rect 9863 2783 16837 2817
<< locali >>
rect 9803 3363 9863 3397
rect 16837 3363 16897 3397
rect 9803 3337 9837 3363
rect 9803 2817 9837 2843
rect 16863 3337 16897 3363
rect 16863 2817 16897 2843
rect 9803 2783 9863 2817
rect 16837 2783 16897 2817
rect 9856 2410 9952 2444
rect 16080 2410 16176 2444
rect 9856 2348 9890 2410
rect 16142 2348 16176 2410
rect 9856 1930 9890 1992
rect 16142 1930 16176 1992
rect 9856 1896 9952 1930
rect 16080 1896 16176 1930
rect 9936 1570 10032 1604
rect 16560 1570 16656 1604
rect 9936 1508 9970 1570
rect 9936 1090 9970 1152
rect 16622 1508 16656 1570
rect 16622 1090 16656 1152
rect 9936 1056 10032 1090
rect 16560 1056 16656 1090
<< viali >>
rect 10420 3397 10540 3420
rect 10420 3363 10540 3397
rect 10420 3360 10540 3363
rect 10280 2300 10440 2340
rect 11060 2300 11220 2340
rect 11300 2300 11460 2340
rect 12080 2300 12240 2340
rect 12340 2300 12500 2340
rect 13120 2300 13280 2340
rect 13380 2300 13540 2340
rect 14140 2300 14300 2340
rect 14400 2300 14560 2340
rect 15180 2300 15340 2340
rect 10020 1980 10180 2020
rect 10540 1980 10700 2020
rect 10800 1980 10960 2020
rect 11560 1980 11720 2020
rect 11820 1980 11980 2020
rect 12600 1980 12760 2020
rect 12860 1980 13020 2020
rect 13640 1980 13800 2020
rect 13880 1980 14040 2020
rect 14660 1980 14820 2020
rect 14920 1980 15080 2020
rect 15440 1980 15600 2020
rect 10160 1090 10500 1100
rect 10160 1056 10500 1090
rect 10160 1040 10500 1056
<< metal1 >>
rect 10400 3440 10600 3620
rect 10170 3360 10180 3440
rect 10240 3420 10700 3440
rect 10240 3380 10420 3420
rect 10240 3360 10250 3380
rect 10408 3360 10420 3380
rect 10540 3380 10700 3420
rect 10540 3360 10552 3380
rect 10690 3360 10700 3380
rect 10760 3360 11200 3440
rect 11260 3380 11580 3440
rect 11640 3380 12220 3440
rect 11260 3360 12220 3380
rect 12280 3360 12740 3440
rect 12800 3360 13240 3440
rect 13300 3360 13640 3440
rect 13700 3360 14140 3440
rect 14200 3360 14660 3440
rect 14720 3360 14800 3440
rect 14860 3360 15440 3440
rect 15500 3360 15960 3440
rect 16020 3360 16480 3440
rect 16540 3360 16550 3440
rect 10408 3354 10552 3360
rect 9960 3180 10180 3260
rect 16520 3180 16740 3260
rect 9920 3000 10180 3180
rect 9960 2900 10180 3000
rect 10240 2980 10250 3180
rect 10410 2980 10420 3180
rect 10480 2980 10490 3180
rect 10690 2980 10700 3180
rect 10760 2980 10770 3180
rect 10930 2980 10940 3180
rect 11000 2980 11010 3180
rect 11190 2980 11200 3180
rect 11260 2980 11270 3180
rect 11450 2980 11460 3180
rect 11520 2980 11530 3180
rect 11570 2980 11580 3180
rect 11640 2980 11650 3180
rect 11810 2980 11820 3180
rect 11880 2980 11890 3180
rect 11950 2980 11960 3180
rect 12020 2980 12030 3180
rect 12210 2980 12220 3180
rect 12280 2980 12290 3180
rect 12470 2980 12480 3180
rect 12540 2980 12550 3180
rect 12710 2980 12720 3180
rect 12780 2980 12790 3180
rect 12970 2980 12980 3180
rect 13040 2980 13050 3180
rect 13230 2980 13240 3180
rect 13300 2980 13310 3180
rect 13370 2980 13380 3180
rect 13440 2980 13450 3180
rect 13630 2980 13640 3180
rect 13700 2980 13710 3180
rect 13890 2980 13900 3180
rect 13960 2980 13970 3180
rect 14130 2980 14140 3180
rect 14200 2980 14210 3180
rect 14390 2980 14400 3180
rect 14460 2980 14470 3180
rect 14650 2980 14660 3180
rect 14720 2980 14730 3180
rect 14790 2980 14800 3180
rect 14860 2980 14870 3180
rect 15050 2980 15130 3180
rect 15170 2980 15180 3180
rect 15240 2980 15250 3180
rect 15430 2980 15440 3180
rect 15500 2980 15510 3180
rect 15670 2980 15680 3180
rect 15740 2980 15750 3180
rect 15950 2980 15960 3180
rect 16020 2980 16030 3180
rect 16210 2980 16220 3180
rect 16280 2980 16290 3180
rect 16470 2980 16480 3180
rect 16540 2980 16780 3180
rect 11840 2940 11880 2980
rect 14910 2940 14990 2980
rect 15060 2940 15120 2980
rect 10240 2900 13240 2940
rect 13440 2920 16460 2940
rect 13440 2900 14840 2920
rect 14830 2860 14840 2900
rect 14900 2900 16460 2920
rect 16520 2900 16740 2980
rect 14900 2860 14910 2900
rect 10400 2720 10420 2800
rect 10480 2780 10500 2800
rect 10930 2780 10940 2800
rect 10480 2720 10940 2780
rect 11000 2780 11010 2800
rect 11450 2780 11460 2800
rect 11000 2720 11340 2780
rect 11400 2720 11460 2780
rect 11520 2780 11530 2800
rect 11950 2780 11960 2800
rect 11520 2720 11960 2780
rect 12020 2780 12030 2800
rect 12470 2780 12480 2800
rect 12020 2720 12480 2780
rect 12540 2780 12550 2800
rect 12970 2780 12980 2800
rect 12540 2720 12980 2780
rect 13040 2720 13050 2800
rect 13350 2720 13360 2800
rect 13420 2780 13430 2800
rect 13870 2780 13880 2800
rect 13420 2720 13880 2780
rect 13940 2780 13950 2800
rect 14390 2780 14400 2800
rect 13940 2720 14400 2780
rect 14460 2780 14470 2800
rect 15170 2780 15180 2800
rect 14460 2720 14720 2780
rect 14780 2720 15180 2780
rect 15240 2780 15250 2800
rect 15670 2780 15680 2800
rect 15240 2720 15680 2780
rect 15740 2780 15750 2800
rect 16210 2780 16220 2800
rect 15740 2720 16220 2780
rect 16280 2720 16290 2800
rect 9760 2660 9960 2720
rect 9760 2600 10300 2660
rect 10360 2600 10370 2660
rect 9760 2520 9960 2600
rect 16720 2580 16920 2600
rect 10450 2500 10460 2560
rect 10520 2500 10820 2560
rect 10880 2500 10980 2560
rect 11040 2500 11480 2560
rect 11540 2500 12000 2560
rect 12060 2500 12520 2560
rect 12580 2500 13040 2560
rect 13100 2500 13540 2560
rect 13600 2500 14060 2560
rect 14120 2500 14580 2560
rect 14640 2500 15100 2560
rect 15160 2500 15170 2560
rect 15230 2520 15240 2580
rect 15300 2520 15720 2580
rect 15240 2500 15720 2520
rect 15780 2500 16920 2580
rect 10170 2380 10180 2440
rect 10240 2380 11220 2440
rect 11280 2380 11820 2440
rect 11880 2380 12260 2440
rect 12320 2380 13280 2440
rect 13340 2380 14320 2440
rect 14380 2380 15360 2440
rect 15420 2380 15440 2440
rect 16720 2400 16920 2500
rect 10268 2340 10452 2346
rect 11048 2340 11232 2346
rect 11288 2340 11472 2346
rect 12068 2340 12252 2346
rect 12328 2340 12512 2346
rect 13108 2340 13292 2346
rect 13368 2340 13552 2346
rect 14128 2340 14312 2346
rect 14388 2340 14572 2346
rect 15168 2340 15352 2346
rect 9980 2260 10220 2340
rect 10268 2300 10280 2340
rect 10440 2300 11060 2340
rect 11220 2300 11300 2340
rect 11460 2300 12080 2340
rect 12240 2300 12340 2340
rect 12500 2300 13120 2340
rect 13280 2300 13380 2340
rect 13540 2300 14140 2340
rect 14300 2300 14400 2340
rect 14560 2300 15180 2340
rect 15340 2300 15352 2340
rect 10268 2294 10452 2300
rect 11048 2294 11232 2300
rect 11288 2294 11472 2300
rect 12068 2294 12252 2300
rect 12328 2294 12512 2300
rect 13108 2294 13292 2300
rect 13368 2294 13552 2300
rect 14128 2294 14312 2300
rect 14388 2294 14572 2300
rect 15168 2294 15240 2300
rect 15230 2280 15240 2294
rect 15300 2294 15352 2300
rect 15300 2280 15310 2294
rect 15400 2260 15640 2340
rect 9980 2060 10180 2260
rect 10240 2060 10250 2260
rect 10450 2060 10460 2260
rect 10520 2060 10530 2260
rect 10690 2060 10700 2260
rect 10760 2060 10770 2260
rect 10970 2060 10980 2260
rect 11040 2060 11050 2260
rect 11210 2060 11220 2260
rect 11280 2060 11290 2260
rect 11470 2060 11480 2260
rect 11540 2060 11550 2260
rect 11730 2060 11740 2260
rect 11800 2060 11810 2260
rect 11990 2060 12000 2260
rect 12060 2060 12070 2260
rect 12250 2060 12260 2260
rect 12320 2060 12330 2260
rect 12510 2060 12520 2260
rect 12580 2060 12590 2260
rect 12770 2070 12780 2250
rect 12840 2070 12850 2250
rect 13030 2060 13040 2260
rect 13100 2060 13110 2260
rect 13270 2060 13280 2260
rect 13340 2060 13350 2260
rect 13530 2060 13540 2260
rect 13600 2060 13610 2260
rect 13790 2060 13800 2260
rect 13860 2060 13870 2260
rect 14050 2060 14060 2260
rect 14120 2060 14130 2260
rect 14310 2060 14320 2260
rect 14380 2060 14390 2260
rect 14570 2060 14580 2260
rect 14640 2060 14650 2260
rect 14830 2250 14900 2260
rect 14830 2060 14840 2250
rect 14900 2060 14910 2250
rect 15400 2240 15680 2260
rect 15090 2060 15100 2240
rect 15160 2060 15170 2240
rect 15350 2060 15360 2240
rect 15420 2080 15680 2240
rect 15420 2060 15640 2080
rect 9980 2020 10220 2060
rect 10290 2020 10300 2040
rect 9980 1980 10020 2020
rect 10180 1980 10220 2020
rect 10280 1980 10300 2020
rect 10360 2020 10370 2040
rect 13670 2026 13750 2040
rect 10528 2020 10712 2026
rect 10788 2020 10972 2026
rect 11548 2020 11732 2026
rect 11808 2020 11992 2026
rect 12588 2020 12772 2026
rect 12848 2020 13032 2026
rect 13628 2020 13812 2026
rect 13868 2020 14052 2026
rect 14648 2020 14832 2026
rect 14908 2020 15092 2026
rect 15400 2020 15640 2060
rect 10360 1980 10540 2020
rect 10700 1980 10800 2020
rect 10960 1980 11560 2020
rect 11720 1980 11820 2020
rect 11980 1980 12600 2020
rect 12760 1980 12860 2020
rect 13020 1980 13640 2020
rect 13800 1980 13880 2020
rect 14040 1980 14660 2020
rect 14820 1980 14920 2020
rect 15080 1980 15340 2020
rect 15400 1980 15440 2020
rect 15600 1980 15640 2020
rect 10008 1974 10192 1980
rect 10528 1974 10712 1980
rect 10788 1974 10972 1980
rect 11548 1974 11732 1980
rect 11808 1974 11992 1980
rect 12588 1974 12772 1980
rect 12848 1974 13032 1980
rect 13628 1974 13812 1980
rect 13868 1974 14052 1980
rect 14648 1974 14832 1980
rect 14908 1974 15092 1980
rect 15428 1974 15612 1980
rect 10680 1880 10700 1940
rect 10760 1880 11740 1940
rect 11800 1880 12780 1940
rect 12840 1880 13800 1940
rect 13860 1880 14840 1940
rect 14900 1880 14910 1940
rect 9760 1780 9960 1840
rect 9760 1720 10300 1780
rect 10360 1720 10370 1780
rect 9760 1640 9960 1720
rect 10930 1680 10940 1740
rect 11000 1680 11340 1740
rect 11400 1680 12000 1740
rect 12060 1680 13020 1740
rect 13080 1680 14060 1740
rect 14120 1680 15080 1740
rect 15140 1680 16120 1740
rect 16180 1680 16190 1740
rect 11470 1560 11480 1620
rect 11540 1560 12520 1620
rect 12580 1560 13540 1620
rect 13600 1560 14560 1620
rect 14620 1560 14720 1620
rect 14780 1560 15600 1620
rect 15660 1560 15720 1620
rect 15780 1560 15790 1620
rect 10080 1420 10260 1500
rect 10060 1260 10300 1420
rect 10080 1160 10260 1260
rect 10290 1240 10300 1260
rect 10360 1280 10370 1420
rect 10820 1380 10920 1420
rect 16220 1400 16440 1500
rect 10360 1240 10440 1280
rect 10550 1240 10560 1380
rect 10620 1240 10630 1380
rect 10810 1240 10820 1380
rect 10880 1260 10920 1380
rect 10880 1240 10890 1260
rect 10950 1240 10960 1400
rect 11020 1300 11030 1400
rect 11020 1240 11080 1300
rect 11210 1240 11220 1400
rect 11280 1240 11290 1400
rect 11470 1240 11480 1400
rect 11540 1240 11550 1400
rect 11730 1240 11740 1400
rect 11800 1240 11810 1400
rect 11990 1240 12000 1400
rect 12060 1240 12070 1400
rect 12250 1240 12260 1400
rect 12320 1240 12330 1400
rect 12510 1240 12520 1400
rect 12580 1240 12590 1400
rect 12750 1240 12760 1400
rect 12820 1240 12830 1400
rect 13010 1240 13020 1400
rect 13080 1240 13090 1400
rect 13270 1240 13280 1400
rect 13340 1240 13350 1400
rect 13530 1240 13540 1400
rect 13600 1240 13610 1400
rect 13790 1240 13800 1400
rect 13860 1240 13870 1400
rect 14050 1240 14060 1400
rect 14120 1240 14130 1400
rect 14310 1240 14320 1400
rect 14380 1240 14390 1400
rect 14550 1240 14560 1400
rect 14620 1240 14650 1400
rect 14810 1240 14820 1400
rect 14880 1240 14910 1400
rect 15070 1240 15080 1400
rect 15140 1240 15150 1400
rect 15330 1240 15340 1400
rect 15400 1240 15410 1400
rect 15590 1240 15600 1400
rect 15660 1240 15670 1400
rect 15850 1240 15860 1400
rect 15920 1240 15930 1400
rect 16110 1240 16120 1400
rect 16180 1260 16440 1400
rect 16180 1240 16190 1260
rect 10340 1200 10440 1240
rect 10980 1200 11080 1240
rect 10340 1180 10800 1200
rect 10360 1160 10800 1180
rect 10980 1160 16080 1200
rect 16220 1160 16440 1260
rect 10148 1100 10512 1106
rect 10148 1080 10160 1100
rect 9760 1040 10160 1080
rect 10500 1080 10512 1100
rect 10500 1040 10560 1080
rect 9760 1020 10560 1040
rect 10620 1020 11220 1080
rect 11280 1020 11740 1080
rect 11800 1020 12260 1080
rect 12320 1020 12760 1080
rect 12820 1020 13280 1080
rect 13340 1020 13800 1080
rect 13860 1020 14320 1080
rect 14380 1020 14820 1080
rect 14880 1020 15340 1080
rect 15400 1020 15860 1080
rect 15920 1020 16190 1080
rect 9760 880 10500 1020
<< via1 >>
rect 10180 3360 10240 3440
rect 10700 3360 10760 3440
rect 11200 3360 11260 3440
rect 11580 3380 11640 3440
rect 12220 3360 12280 3440
rect 12740 3360 12800 3440
rect 13240 3360 13300 3440
rect 13640 3360 13700 3440
rect 14140 3360 14200 3440
rect 14660 3360 14720 3440
rect 14800 3360 14860 3440
rect 15440 3360 15500 3440
rect 15960 3360 16020 3440
rect 16480 3360 16540 3440
rect 10180 2980 10240 3180
rect 10420 2980 10480 3180
rect 10700 2980 10760 3180
rect 10940 2980 11000 3180
rect 11200 2980 11260 3180
rect 11460 2980 11520 3180
rect 11580 2980 11640 3180
rect 11820 2980 11880 3180
rect 11960 2980 12020 3180
rect 12220 2980 12280 3180
rect 12480 2980 12540 3180
rect 12720 2980 12780 3180
rect 12980 2980 13040 3180
rect 13240 2980 13300 3180
rect 13380 2980 13440 3180
rect 13640 2980 13700 3180
rect 13900 2980 13960 3180
rect 14140 2980 14200 3180
rect 14400 2980 14460 3180
rect 14660 2980 14720 3180
rect 14800 2980 14860 3180
rect 15180 2980 15240 3180
rect 15440 2980 15500 3180
rect 15680 2980 15740 3180
rect 15960 2980 16020 3180
rect 16220 2980 16280 3180
rect 16480 2980 16540 3180
rect 14840 2860 14900 2920
rect 10420 2720 10480 2800
rect 10940 2720 11000 2800
rect 11340 2720 11400 2780
rect 11460 2720 11520 2800
rect 11960 2720 12020 2800
rect 12480 2720 12540 2800
rect 12980 2720 13040 2800
rect 13360 2720 13420 2800
rect 13880 2720 13940 2800
rect 14400 2720 14460 2800
rect 14720 2720 14780 2780
rect 15180 2720 15240 2800
rect 15680 2720 15740 2800
rect 16220 2720 16280 2800
rect 10300 2600 10360 2660
rect 10460 2500 10520 2560
rect 10820 2500 10880 2560
rect 10980 2500 11040 2560
rect 11480 2500 11540 2560
rect 12000 2500 12060 2560
rect 12520 2500 12580 2560
rect 13040 2500 13100 2560
rect 13540 2500 13600 2560
rect 14060 2500 14120 2560
rect 14580 2500 14640 2560
rect 15100 2500 15160 2560
rect 15240 2520 15300 2580
rect 15720 2500 15780 2580
rect 10180 2380 10240 2440
rect 11220 2380 11280 2440
rect 11820 2380 11880 2440
rect 12260 2380 12320 2440
rect 13280 2380 13340 2440
rect 14320 2380 14380 2440
rect 15360 2380 15420 2440
rect 15240 2300 15300 2340
rect 15240 2280 15300 2300
rect 10180 2060 10240 2260
rect 10460 2060 10520 2260
rect 10700 2060 10760 2260
rect 10980 2060 11040 2260
rect 11220 2060 11280 2260
rect 11480 2060 11540 2260
rect 11740 2060 11800 2260
rect 12000 2060 12060 2260
rect 12260 2060 12320 2260
rect 12520 2060 12580 2260
rect 12780 2070 12840 2250
rect 13040 2060 13100 2260
rect 13280 2060 13340 2260
rect 13540 2060 13600 2260
rect 13800 2060 13860 2260
rect 14060 2060 14120 2260
rect 14320 2060 14380 2260
rect 14580 2060 14640 2260
rect 14840 2060 14900 2250
rect 15100 2060 15160 2240
rect 15360 2060 15420 2240
rect 10300 1980 10360 2040
rect 10700 1880 10760 1940
rect 11740 1880 11800 1940
rect 12780 1880 12840 1940
rect 13800 1880 13860 1940
rect 14840 1880 14900 1940
rect 10300 1720 10360 1780
rect 10940 1680 11000 1740
rect 11340 1680 11400 1740
rect 12000 1680 12060 1740
rect 13020 1680 13080 1740
rect 14060 1680 14120 1740
rect 15080 1680 15140 1740
rect 16120 1680 16180 1740
rect 11480 1560 11540 1620
rect 12520 1560 12580 1620
rect 13540 1560 13600 1620
rect 14560 1560 14620 1620
rect 14720 1560 14780 1620
rect 15600 1560 15660 1620
rect 15720 1560 15780 1620
rect 10300 1240 10360 1420
rect 10560 1240 10620 1380
rect 10820 1240 10880 1380
rect 10960 1240 11020 1400
rect 11220 1240 11280 1400
rect 11480 1240 11540 1400
rect 11740 1240 11800 1400
rect 12000 1240 12060 1400
rect 12260 1240 12320 1400
rect 12520 1240 12580 1400
rect 12760 1240 12820 1400
rect 13020 1240 13080 1400
rect 13280 1240 13340 1400
rect 13540 1240 13600 1400
rect 13800 1240 13860 1400
rect 14060 1240 14120 1400
rect 14320 1240 14380 1400
rect 14560 1240 14620 1400
rect 14820 1240 14880 1400
rect 15080 1240 15140 1400
rect 15340 1240 15400 1400
rect 15600 1240 15660 1400
rect 15860 1240 15920 1400
rect 16120 1240 16180 1400
rect 10560 1020 10620 1080
rect 11220 1020 11280 1080
rect 11740 1020 11800 1080
rect 12260 1020 12320 1080
rect 12760 1020 12820 1080
rect 13280 1020 13340 1080
rect 13800 1020 13860 1080
rect 14320 1020 14380 1080
rect 14820 1020 14880 1080
rect 15340 1020 15400 1080
rect 15860 1020 15920 1080
<< metal2 >>
rect 10180 3440 10240 3450
rect 10180 3180 10240 3360
rect 10700 3440 10760 3450
rect 10180 2970 10240 2980
rect 10420 3180 10480 3190
rect 10420 2800 10480 2980
rect 10700 3180 10760 3360
rect 11200 3440 11260 3450
rect 10700 2970 10760 2980
rect 10940 3180 11000 3190
rect 10420 2710 10480 2720
rect 10940 2800 11000 2980
rect 11200 3180 11260 3360
rect 11580 3440 11640 3450
rect 11200 2970 11260 2980
rect 11460 3180 11520 3190
rect 11460 2800 11520 2980
rect 11580 3180 11640 3380
rect 12220 3440 12280 3450
rect 11580 2970 11640 2980
rect 11820 3180 11880 3190
rect 10940 2710 11000 2720
rect 11340 2780 11400 2800
rect 10300 2660 10360 2670
rect 10180 2440 10240 2460
rect 10180 2260 10240 2380
rect 10180 2050 10240 2060
rect 10300 2040 10360 2600
rect 10460 2560 10520 2570
rect 10460 2260 10520 2500
rect 10820 2560 10880 2570
rect 10460 2050 10520 2060
rect 10700 2260 10760 2270
rect 10300 1970 10360 1980
rect 10700 1940 10760 2060
rect 10700 1870 10760 1880
rect 10300 1780 10360 1790
rect 10300 1420 10360 1720
rect 10300 1230 10360 1240
rect 10560 1380 10620 1390
rect 10560 1080 10620 1240
rect 10820 1380 10880 2500
rect 10980 2560 11040 2570
rect 10980 2260 11040 2500
rect 10980 2050 11040 2060
rect 11220 2440 11280 2450
rect 11220 2260 11280 2380
rect 11220 2050 11280 2060
rect 10820 1230 10880 1240
rect 10940 1740 11000 1750
rect 10940 1410 11000 1680
rect 11340 1740 11400 2720
rect 11460 2710 11520 2720
rect 11480 2560 11540 2570
rect 11480 2260 11540 2500
rect 11820 2440 11880 2980
rect 11960 3180 12020 3190
rect 11960 2800 12020 2980
rect 12220 3180 12280 3360
rect 12740 3440 12800 3450
rect 12740 3190 12800 3360
rect 13240 3440 13300 3450
rect 12220 2970 12280 2980
rect 12480 3180 12540 3190
rect 11960 2710 12020 2720
rect 12480 2800 12540 2980
rect 12720 3180 12800 3190
rect 12780 2980 12800 3180
rect 12980 3180 13040 3190
rect 12720 2970 12780 2980
rect 12480 2710 12540 2720
rect 12980 2800 13040 2980
rect 13240 3180 13300 3360
rect 13640 3440 13700 3450
rect 13380 3180 13440 3190
rect 13240 2970 13300 2980
rect 13360 2980 13380 3180
rect 13360 2970 13440 2980
rect 13640 3180 13700 3360
rect 14140 3440 14200 3450
rect 13900 3180 13960 3190
rect 13640 2970 13700 2980
rect 13880 2980 13900 3180
rect 13880 2970 13960 2980
rect 14140 3180 14200 3360
rect 14660 3440 14720 3450
rect 14140 2970 14200 2980
rect 14400 3180 14460 3190
rect 12980 2710 13040 2720
rect 13360 2800 13420 2970
rect 13360 2710 13420 2720
rect 13880 2800 13940 2970
rect 13880 2710 13940 2720
rect 14400 2800 14460 2980
rect 14660 3180 14720 3360
rect 14660 2970 14720 2980
rect 14800 3440 14860 3450
rect 14800 3180 14860 3360
rect 15440 3440 15500 3450
rect 14800 2970 14860 2980
rect 15180 3180 15240 3190
rect 14840 2920 14900 2940
rect 14400 2700 14460 2720
rect 14720 2780 14780 2790
rect 11820 2370 11880 2380
rect 12000 2560 12060 2570
rect 11480 2050 11540 2060
rect 11740 2260 11800 2270
rect 11740 1940 11800 2060
rect 12000 2260 12060 2500
rect 12520 2560 12580 2570
rect 12000 2050 12060 2060
rect 12260 2440 12320 2450
rect 12260 2260 12320 2380
rect 12260 2050 12320 2060
rect 12520 2260 12580 2500
rect 13040 2560 13100 2570
rect 13040 2260 13100 2500
rect 13540 2560 13600 2570
rect 12520 2050 12580 2060
rect 12780 2250 12840 2260
rect 11740 1870 11800 1880
rect 12780 1940 12840 2070
rect 13040 2050 13100 2060
rect 13280 2440 13340 2450
rect 13280 2260 13340 2380
rect 13280 2050 13340 2060
rect 13540 2260 13600 2500
rect 14060 2560 14120 2570
rect 13540 2050 13600 2060
rect 13800 2260 13860 2270
rect 12780 1870 12840 1880
rect 13800 1940 13860 2060
rect 14060 2260 14120 2500
rect 14580 2560 14640 2570
rect 14060 2050 14120 2060
rect 14320 2440 14380 2450
rect 14320 2260 14380 2380
rect 14320 2050 14380 2060
rect 14580 2260 14640 2500
rect 14580 2050 14640 2060
rect 13800 1870 13860 1880
rect 11340 1670 11400 1680
rect 12000 1740 12060 1750
rect 11480 1620 11540 1630
rect 10940 1400 11020 1410
rect 10940 1240 10960 1400
rect 10940 1230 11020 1240
rect 11220 1400 11280 1410
rect 10560 1010 10620 1020
rect 10940 700 11000 1230
rect 11220 1080 11280 1240
rect 11480 1400 11540 1560
rect 11480 1230 11540 1240
rect 11740 1400 11800 1410
rect 11220 1010 11280 1020
rect 11740 1080 11800 1240
rect 12000 1400 12060 1680
rect 13020 1740 13080 1750
rect 12520 1620 12580 1630
rect 12000 1230 12060 1240
rect 12260 1400 12320 1410
rect 11740 1010 11800 1020
rect 12260 1080 12320 1240
rect 12520 1400 12580 1560
rect 12520 1230 12580 1240
rect 12760 1400 12820 1410
rect 12260 1010 12320 1020
rect 12760 1080 12820 1240
rect 13020 1400 13080 1680
rect 14060 1740 14120 1750
rect 13540 1620 13600 1630
rect 13020 1220 13080 1240
rect 13280 1400 13340 1410
rect 12760 1010 12820 1020
rect 13280 1080 13340 1240
rect 13540 1400 13600 1560
rect 13540 1220 13600 1240
rect 13800 1400 13860 1410
rect 13280 1010 13340 1020
rect 13800 1080 13860 1240
rect 14060 1400 14120 1680
rect 14560 1620 14620 1630
rect 14060 1220 14120 1240
rect 14320 1400 14380 1410
rect 13800 1010 13860 1020
rect 14320 1080 14380 1240
rect 14560 1400 14620 1560
rect 14720 1620 14780 2720
rect 14840 2260 14900 2860
rect 15180 2800 15240 2980
rect 15440 3180 15500 3360
rect 15960 3440 16020 3450
rect 15440 2970 15500 2980
rect 15680 3180 15740 3190
rect 15180 2710 15240 2720
rect 15680 2800 15740 2980
rect 15960 3180 16020 3360
rect 16480 3440 16540 3450
rect 15960 2970 16020 2980
rect 16220 3180 16280 3190
rect 15680 2710 15740 2720
rect 16220 2800 16280 2980
rect 16480 3180 16540 3360
rect 16480 2970 16540 2980
rect 16220 2710 16280 2720
rect 15240 2580 15300 2590
rect 14830 2250 14900 2260
rect 14830 2060 14840 2250
rect 14840 1940 14900 2060
rect 15100 2560 15160 2570
rect 15100 2240 15160 2500
rect 15240 2340 15300 2520
rect 15720 2580 15780 2590
rect 15240 2270 15300 2280
rect 15360 2440 15420 2450
rect 15100 2050 15160 2060
rect 15360 2240 15420 2380
rect 15360 2050 15420 2060
rect 14840 1870 14900 1880
rect 14720 1540 14780 1560
rect 15080 1740 15140 1750
rect 14560 1220 14620 1240
rect 14820 1400 14880 1410
rect 14320 1010 14380 1020
rect 14820 1080 14880 1240
rect 15080 1400 15140 1680
rect 15600 1620 15660 1630
rect 15080 1220 15140 1240
rect 15340 1400 15400 1410
rect 14820 1010 14880 1020
rect 15340 1080 15400 1240
rect 15600 1400 15660 1560
rect 15600 1220 15660 1240
rect 15720 1620 15780 2500
rect 15340 1010 15400 1020
rect 15720 960 15780 1560
rect 16120 1740 16180 1750
rect 15860 1400 15920 1410
rect 15860 1080 15920 1240
rect 16120 1400 16180 1680
rect 16120 1220 16180 1240
rect 15860 1010 15920 1020
rect 15720 870 15780 880
rect 10940 610 11000 620
<< via2 >>
rect 15720 880 15780 960
rect 10940 620 11000 700
<< metal3 >>
rect 15710 960 15790 965
rect 15710 940 15720 960
rect 15680 880 15720 940
rect 15780 940 15790 960
rect 15780 920 16320 940
rect 15780 880 16080 920
rect 15680 860 16080 880
rect 16070 720 16080 860
rect 16380 720 16390 920
rect 10930 700 11010 705
rect 10130 620 10140 700
rect 10260 620 10940 700
rect 11000 620 11010 700
rect 10930 615 11010 620
<< via3 >>
rect 16080 720 16380 920
rect 10140 620 10260 700
<< metal4 >>
rect 10139 700 10261 701
rect 10139 620 10140 700
rect 10260 620 10261 700
rect 10139 619 10261 620
rect 10160 280 10240 619
<< via4 >>
rect 16040 920 16400 940
rect 16040 720 16080 920
rect 16080 720 16380 920
rect 16380 720 16400 920
rect 16040 660 16400 720
<< metal5 >>
rect 16016 940 16424 964
rect 16016 660 16040 940
rect 16400 660 16424 940
rect 16016 636 16424 660
rect 16060 60 16400 636
use sky130_fd_pr__cap_mim_m3_2_26U9NK  sky130_fd_pr__cap_mim_m3_2_26U9NK_0
timestamp 1700064502
transform -1 0 13431 0 -1 -1279
box -3349 -1581 3371 1581
use sky130_fd_pr__nfet_01v8_HBAYNJ  sky130_fd_pr__nfet_01v8_HBAYNJ_0
timestamp 1700066397
transform 1 0 12813 0 1 2162
box -2867 -188 2867 188
use sky130_fd_pr__nfet_01v8_XWAA4X  sky130_fd_pr__nfet_01v8_XWAA4X_0
timestamp 1700070217
transform 1 0 10456 0 1 1328
box -416 -188 416 188
use sky130_fd_pr__pfet_01v8_3H5TVM  sky130_fd_pr__pfet_01v8_3H5TVM_0
timestamp 1700009976
transform 1 0 11734 0 1 3080
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_3H5TVM  sky130_fd_pr__pfet_01v8_3H5TVM_1
timestamp 1700009976
transform 1 0 14954 0 1 3080
box -194 -200 194 200
use sky130_fd_pr__pfet_01v8_3HMWVM  sky130_fd_pr__pfet_01v8_3HMWVM_0
timestamp 1700012548
transform 1 0 12630 0 1 3080
box -710 -200 710 200
use sky130_fd_pr__pfet_01v8_3HMWVM  sky130_fd_pr__pfet_01v8_3HMWVM_3
timestamp 1700012548
transform 1 0 14050 0 1 3080
box -710 -200 710 200
use sky130_fd_pr__pfet_01v8_3HZSVM  sky130_fd_pr__pfet_01v8_3HZSVM_0
timestamp 1700012548
transform 1 0 10719 0 1 3080
box -839 -200 839 200
use sky130_fd_pr__pfet_01v8_3HZSVM  sky130_fd_pr__pfet_01v8_3HZSVM_1
timestamp 1700012548
transform 1 0 15979 0 1 3080
box -839 -200 839 200
use sky130_fd_pr__nfet_01v8_P8B44K  XM9
timestamp 1700063261
transform 1 0 13698 0 1 1328
box -2738 -188 2738 188
<< labels >>
flabel metal1 10400 3420 10600 3620 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal2 11360 1800 11380 1820 0 FreeSans 800 0 0 0 d
flabel metal1 16720 2400 16920 2600 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 9760 2520 9960 2720 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal2 11820 2660 11840 2660 0 FreeSans 800 0 0 0 a
flabel metal2 10840 1800 10860 1820 0 FreeSans 800 0 0 0 c
flabel metal2 14860 2640 14860 2640 0 FreeSans 800 0 0 0 b
flabel metal1 9760 1640 9960 1840 0 FreeSans 256 0 0 0 ib
port 1 nsew
flabel metal1 9760 880 9960 1080 0 FreeSans 256 0 0 0 gnd
port 6 nsew
<< end >>
