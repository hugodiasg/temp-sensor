magic
tech sky130A
magscale 1 2
timestamp 1646183319
<< metal4 >>
rect -2481 7265 2481 7306
rect -2481 2543 2225 7265
rect 2461 2543 2481 7265
rect -2481 2502 2481 2543
rect -2481 2361 2481 2402
rect -2481 -2361 2225 2361
rect 2461 -2361 2481 2361
rect -2481 -2402 2481 -2361
rect -2481 -2543 2481 -2502
rect -2481 -7265 2225 -2543
rect 2461 -7265 2481 -2543
rect -2481 -7306 2481 -7265
<< via4 >>
rect 2225 2543 2461 7265
rect 2225 -2361 2461 2361
rect 2225 -7265 2461 -2543
<< mimcap2 >>
rect -2381 7166 2223 7206
rect -2381 2642 -1889 7166
rect 1731 2642 2223 7166
rect -2381 2602 2223 2642
rect -2381 2262 2223 2302
rect -2381 -2262 -1889 2262
rect 1731 -2262 2223 2262
rect -2381 -2302 2223 -2262
rect -2381 -2642 2223 -2602
rect -2381 -7166 -1889 -2642
rect 1731 -7166 2223 -2642
rect -2381 -7206 2223 -7166
<< mimcap2contact >>
rect -1889 2642 1731 7166
rect -1889 -2262 1731 2262
rect -1889 -7166 1731 -2642
<< metal5 >>
rect -239 7190 81 7356
rect 2183 7265 2503 7356
rect -1913 7166 1755 7190
rect -1913 2642 -1889 7166
rect 1731 2642 1755 7166
rect -1913 2618 1755 2642
rect -239 2286 81 2618
rect 2183 2543 2225 7265
rect 2461 2543 2503 7265
rect 2183 2361 2503 2543
rect -1913 2262 1755 2286
rect -1913 -2262 -1889 2262
rect 1731 -2262 1755 2262
rect -1913 -2286 1755 -2262
rect -239 -2618 81 -2286
rect 2183 -2361 2225 2361
rect 2461 -2361 2503 2361
rect 2183 -2543 2503 -2361
rect -1913 -2642 1755 -2618
rect -1913 -7166 -1889 -2642
rect 1731 -7166 1755 -2642
rect -1913 -7190 1755 -7166
rect -239 -7356 81 -7190
rect 2183 -7265 2225 -2543
rect 2461 -7265 2503 -2543
rect 2183 -7356 2503 -7265
<< properties >>
string FIXED_BBOX -2481 2502 2323 7306
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.016 l 23.016 val 1.076k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
