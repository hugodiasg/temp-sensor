magic
tech sky130A
magscale 1 2
timestamp 1668746776
<< nwell >>
rect -5700 2120 -5108 3758
rect -3140 2120 -2548 3758
rect -540 2100 52 3738
rect 5720 2880 6312 3518
rect 5720 1960 6312 2598
rect -5700 780 -5108 1818
rect -3140 760 -2548 1798
rect -540 740 60 1780
<< pwell >>
rect 1280 1140 1872 1760
rect 7600 1140 8192 1760
rect -5700 60 -5108 680
rect -3140 60 -2548 680
rect -520 40 40 660
rect 360 260 952 880
rect 7600 260 8192 880
<< nmos >>
rect 1476 1350 1676 1550
rect 7796 1350 7996 1550
rect -5504 270 -5304 470
rect -2944 270 -2744 470
rect -344 250 -144 450
rect 556 470 756 670
rect 7796 470 7996 670
<< pmos >>
rect -5504 2339 -5304 3539
rect -2944 2339 -2744 3539
rect -344 2319 -144 3519
rect 5916 3099 6116 3299
rect 5916 2179 6116 2379
rect -5504 999 -5304 1599
rect -2944 979 -2744 1579
rect -344 959 -144 1559
<< ndiff >>
rect 1418 1538 1476 1550
rect 1418 1362 1430 1538
rect 1464 1362 1476 1538
rect 1418 1350 1476 1362
rect 1676 1538 1734 1550
rect 1676 1362 1688 1538
rect 1722 1362 1734 1538
rect 1676 1350 1734 1362
rect 7738 1538 7796 1550
rect 7738 1362 7750 1538
rect 7784 1362 7796 1538
rect 7738 1350 7796 1362
rect 7996 1538 8054 1550
rect 7996 1362 8008 1538
rect 8042 1362 8054 1538
rect 7996 1350 8054 1362
rect -5562 458 -5504 470
rect -5562 282 -5550 458
rect -5516 282 -5504 458
rect -5562 270 -5504 282
rect -5304 458 -5246 470
rect -5304 282 -5292 458
rect -5258 282 -5246 458
rect -5304 270 -5246 282
rect -3002 458 -2944 470
rect -3002 282 -2990 458
rect -2956 282 -2944 458
rect -3002 270 -2944 282
rect -2744 458 -2686 470
rect -2744 282 -2732 458
rect -2698 282 -2686 458
rect -2744 270 -2686 282
rect -402 438 -344 450
rect -402 262 -390 438
rect -356 262 -344 438
rect -402 250 -344 262
rect -144 438 -86 450
rect -144 262 -132 438
rect -98 262 -86 438
rect -144 250 -86 262
rect 498 658 556 670
rect 498 482 510 658
rect 544 482 556 658
rect 498 470 556 482
rect 756 658 814 670
rect 756 482 768 658
rect 802 482 814 658
rect 756 470 814 482
rect 7738 658 7796 670
rect 7738 482 7750 658
rect 7784 482 7796 658
rect 7738 470 7796 482
rect 7996 658 8054 670
rect 7996 482 8008 658
rect 8042 482 8054 658
rect 7996 470 8054 482
<< pdiff >>
rect -5562 3527 -5504 3539
rect -5562 2351 -5550 3527
rect -5516 2351 -5504 3527
rect -5562 2339 -5504 2351
rect -5304 3527 -5246 3539
rect -5304 2351 -5292 3527
rect -5258 2351 -5246 3527
rect -5304 2339 -5246 2351
rect -3002 3527 -2944 3539
rect -3002 2351 -2990 3527
rect -2956 2351 -2944 3527
rect -3002 2339 -2944 2351
rect -2744 3527 -2686 3539
rect -2744 2351 -2732 3527
rect -2698 2351 -2686 3527
rect -2744 2339 -2686 2351
rect -402 3507 -344 3519
rect -402 2331 -390 3507
rect -356 2331 -344 3507
rect -402 2319 -344 2331
rect -144 3507 -86 3519
rect -144 2331 -132 3507
rect -98 2331 -86 3507
rect -144 2319 -86 2331
rect 5858 3287 5916 3299
rect 5858 3111 5870 3287
rect 5904 3111 5916 3287
rect 5858 3099 5916 3111
rect 6116 3287 6174 3299
rect 6116 3111 6128 3287
rect 6162 3111 6174 3287
rect 6116 3099 6174 3111
rect 5858 2367 5916 2379
rect 5858 2191 5870 2367
rect 5904 2191 5916 2367
rect 5858 2179 5916 2191
rect 6116 2367 6174 2379
rect 6116 2191 6128 2367
rect 6162 2191 6174 2367
rect 6116 2179 6174 2191
rect -5562 1587 -5504 1599
rect -5562 1011 -5550 1587
rect -5516 1011 -5504 1587
rect -5562 999 -5504 1011
rect -5304 1587 -5246 1599
rect -5304 1011 -5292 1587
rect -5258 1011 -5246 1587
rect -5304 999 -5246 1011
rect -3002 1567 -2944 1579
rect -3002 991 -2990 1567
rect -2956 991 -2944 1567
rect -3002 979 -2944 991
rect -2744 1567 -2686 1579
rect -2744 991 -2732 1567
rect -2698 991 -2686 1567
rect -2744 979 -2686 991
rect -402 1547 -344 1559
rect -402 971 -390 1547
rect -356 971 -344 1547
rect -402 959 -344 971
rect -144 1547 -86 1559
rect -144 971 -132 1547
rect -98 971 -86 1547
rect -144 959 -86 971
<< ndiffc >>
rect 1430 1362 1464 1538
rect 1688 1362 1722 1538
rect 7750 1362 7784 1538
rect 8008 1362 8042 1538
rect -5550 282 -5516 458
rect -5292 282 -5258 458
rect -2990 282 -2956 458
rect -2732 282 -2698 458
rect -390 262 -356 438
rect -132 262 -98 438
rect 510 482 544 658
rect 768 482 802 658
rect 7750 482 7784 658
rect 8008 482 8042 658
<< pdiffc >>
rect -5550 2351 -5516 3527
rect -5292 2351 -5258 3527
rect -2990 2351 -2956 3527
rect -2732 2351 -2698 3527
rect -390 2331 -356 3507
rect -132 2331 -98 3507
rect 5870 3111 5904 3287
rect 6128 3111 6162 3287
rect 5870 2191 5904 2367
rect 6128 2191 6162 2367
rect -5550 1011 -5516 1587
rect -5292 1011 -5258 1587
rect -2990 991 -2956 1567
rect -2732 991 -2698 1567
rect -390 971 -356 1547
rect -132 971 -98 1547
<< psubdiff >>
rect 1316 1690 1412 1724
rect 1740 1690 1836 1724
rect 1316 1628 1350 1690
rect 1802 1628 1836 1690
rect 1316 1210 1350 1272
rect 1802 1210 1836 1272
rect 1316 1176 1412 1210
rect 1740 1176 1836 1210
rect 7636 1690 7732 1724
rect 8060 1690 8156 1724
rect 7636 1628 7670 1690
rect 8122 1628 8156 1690
rect 7636 1210 7670 1272
rect 8122 1210 8156 1272
rect 7636 1176 7732 1210
rect 8060 1176 8156 1210
rect 396 810 492 844
rect 820 810 916 844
rect 396 748 430 810
rect -5664 610 -5568 644
rect -5240 610 -5144 644
rect -5664 548 -5630 610
rect -5178 548 -5144 610
rect -5664 130 -5630 192
rect -5178 130 -5144 192
rect -5664 96 -5568 130
rect -5240 96 -5144 130
rect -3104 610 -3008 644
rect -2680 610 -2584 644
rect -3104 548 -3070 610
rect -2618 548 -2584 610
rect -3104 130 -3070 192
rect -2618 130 -2584 192
rect -3104 96 -3008 130
rect -2680 96 -2584 130
rect -504 590 -408 624
rect -80 590 16 624
rect -504 528 -470 590
rect -18 528 16 590
rect -504 110 -470 172
rect 882 748 916 810
rect 396 330 430 392
rect 882 330 916 392
rect 396 296 492 330
rect 820 296 916 330
rect 7636 810 7732 844
rect 8060 810 8156 844
rect 7636 748 7670 810
rect 8122 748 8156 810
rect 7636 330 7670 392
rect 8122 330 8156 392
rect 7636 296 7732 330
rect 8060 296 8156 330
rect -18 110 16 172
rect -504 76 -408 110
rect -80 76 16 110
<< nsubdiff >>
rect -5664 3688 -5568 3722
rect -5240 3688 -5144 3722
rect -5664 3626 -5630 3688
rect -5178 3626 -5144 3688
rect -5664 2190 -5630 2252
rect -5178 2190 -5144 2252
rect -5664 2156 -5568 2190
rect -5240 2156 -5144 2190
rect -3104 3688 -3008 3722
rect -2680 3688 -2584 3722
rect -3104 3626 -3070 3688
rect -2618 3626 -2584 3688
rect -3104 2190 -3070 2252
rect -2618 2190 -2584 2252
rect -3104 2156 -3008 2190
rect -2680 2156 -2584 2190
rect -504 3668 -408 3702
rect -80 3668 16 3702
rect -504 3606 -470 3668
rect -18 3606 16 3668
rect -504 2170 -470 2232
rect 5756 3448 5852 3482
rect 6180 3448 6276 3482
rect 5756 3386 5790 3448
rect 6242 3386 6276 3448
rect 5756 2950 5790 3012
rect 6242 2950 6276 3012
rect 5756 2916 5852 2950
rect 6180 2916 6276 2950
rect -18 2170 16 2232
rect -504 2136 -408 2170
rect -80 2136 16 2170
rect 5756 2528 5852 2562
rect 6180 2528 6276 2562
rect 5756 2466 5790 2528
rect 6242 2466 6276 2528
rect 5756 2030 5790 2092
rect 6242 2030 6276 2092
rect 5756 1996 5852 2030
rect 6180 1996 6276 2030
rect -5664 1748 -5568 1782
rect -5240 1748 -5144 1782
rect -5664 1686 -5630 1748
rect -5178 1686 -5144 1748
rect -5664 850 -5630 912
rect -5178 850 -5144 912
rect -5664 816 -5568 850
rect -5240 816 -5144 850
rect -3104 1728 -3008 1762
rect -2680 1728 -2584 1762
rect -3104 1666 -3070 1728
rect -2618 1666 -2584 1728
rect -3104 830 -3070 892
rect -2618 830 -2584 892
rect -3104 796 -3008 830
rect -2680 796 -2584 830
rect -504 1708 -408 1742
rect -80 1708 16 1742
rect -504 1646 -470 1708
rect -18 1646 16 1708
rect -504 810 -470 872
rect -18 810 16 872
rect -504 776 -408 810
rect -80 776 16 810
<< psubdiffcont >>
rect 1412 1690 1740 1724
rect 1316 1272 1350 1628
rect 1802 1272 1836 1628
rect 1412 1176 1740 1210
rect 7732 1690 8060 1724
rect 7636 1272 7670 1628
rect 8122 1272 8156 1628
rect 7732 1176 8060 1210
rect 492 810 820 844
rect -5568 610 -5240 644
rect -5664 192 -5630 548
rect -5178 192 -5144 548
rect -5568 96 -5240 130
rect -3008 610 -2680 644
rect -3104 192 -3070 548
rect -2618 192 -2584 548
rect -3008 96 -2680 130
rect -408 590 -80 624
rect -504 172 -470 528
rect -18 172 16 528
rect 396 392 430 748
rect 882 392 916 748
rect 492 296 820 330
rect 7732 810 8060 844
rect 7636 392 7670 748
rect 8122 392 8156 748
rect 7732 296 8060 330
rect -408 76 -80 110
<< nsubdiffcont >>
rect -5568 3688 -5240 3722
rect -5664 2252 -5630 3626
rect -5178 2252 -5144 3626
rect -5568 2156 -5240 2190
rect -3008 3688 -2680 3722
rect -3104 2252 -3070 3626
rect -2618 2252 -2584 3626
rect -3008 2156 -2680 2190
rect -408 3668 -80 3702
rect -504 2232 -470 3606
rect -18 2232 16 3606
rect 5852 3448 6180 3482
rect 5756 3012 5790 3386
rect 6242 3012 6276 3386
rect 5852 2916 6180 2950
rect -408 2136 -80 2170
rect 5852 2528 6180 2562
rect 5756 2092 5790 2466
rect 6242 2092 6276 2466
rect 5852 1996 6180 2030
rect -5568 1748 -5240 1782
rect -5664 912 -5630 1686
rect -5178 912 -5144 1686
rect -5568 816 -5240 850
rect -3008 1728 -2680 1762
rect -3104 892 -3070 1666
rect -2618 892 -2584 1666
rect -3008 796 -2680 830
rect -408 1708 -80 1742
rect -504 872 -470 1646
rect -18 872 16 1646
rect -408 776 -80 810
<< poly >>
rect -5504 3620 -5304 3636
rect -5504 3586 -5488 3620
rect -5320 3586 -5304 3620
rect -5504 3539 -5304 3586
rect -5504 2292 -5304 2339
rect -5504 2258 -5488 2292
rect -5320 2258 -5304 2292
rect -5504 2242 -5304 2258
rect -2944 3620 -2744 3636
rect -2944 3586 -2928 3620
rect -2760 3586 -2744 3620
rect -2944 3539 -2744 3586
rect -2944 2292 -2744 2339
rect -2944 2258 -2928 2292
rect -2760 2258 -2744 2292
rect -2944 2242 -2744 2258
rect -344 3600 -144 3616
rect -344 3566 -328 3600
rect -160 3566 -144 3600
rect -344 3519 -144 3566
rect -344 2272 -144 2319
rect -344 2238 -328 2272
rect -160 2238 -144 2272
rect -344 2222 -144 2238
rect 5916 3380 6116 3396
rect 5916 3346 5932 3380
rect 6100 3346 6116 3380
rect 5916 3299 6116 3346
rect 5916 3052 6116 3099
rect 5916 3018 5932 3052
rect 6100 3018 6116 3052
rect 5916 3002 6116 3018
rect 5916 2460 6116 2476
rect 5916 2426 5932 2460
rect 6100 2426 6116 2460
rect 5916 2379 6116 2426
rect 5916 2132 6116 2179
rect 5916 2098 5932 2132
rect 6100 2098 6116 2132
rect 5916 2082 6116 2098
rect -5504 1680 -5304 1696
rect -5504 1646 -5488 1680
rect -5320 1646 -5304 1680
rect -5504 1599 -5304 1646
rect -5504 952 -5304 999
rect -5504 918 -5488 952
rect -5320 918 -5304 952
rect -5504 902 -5304 918
rect -2944 1660 -2744 1676
rect -2944 1626 -2928 1660
rect -2760 1626 -2744 1660
rect -2944 1579 -2744 1626
rect -2944 932 -2744 979
rect -2944 898 -2928 932
rect -2760 898 -2744 932
rect -2944 882 -2744 898
rect -344 1640 -144 1656
rect -344 1606 -328 1640
rect -160 1606 -144 1640
rect -344 1559 -144 1606
rect -344 912 -144 959
rect -344 878 -328 912
rect -160 878 -144 912
rect -344 862 -144 878
rect 1476 1622 1676 1638
rect 1476 1588 1492 1622
rect 1660 1588 1676 1622
rect 1476 1550 1676 1588
rect 1476 1312 1676 1350
rect 1476 1278 1492 1312
rect 1660 1278 1676 1312
rect 1476 1262 1676 1278
rect 7796 1622 7996 1638
rect 7796 1588 7812 1622
rect 7980 1588 7996 1622
rect 7796 1550 7996 1588
rect 7796 1312 7996 1350
rect 7796 1278 7812 1312
rect 7980 1278 7996 1312
rect 7796 1262 7996 1278
rect -5504 542 -5304 558
rect -5504 508 -5488 542
rect -5320 508 -5304 542
rect -5504 470 -5304 508
rect -5504 232 -5304 270
rect -5504 198 -5488 232
rect -5320 198 -5304 232
rect -5504 182 -5304 198
rect -2944 542 -2744 558
rect -2944 508 -2928 542
rect -2760 508 -2744 542
rect -2944 470 -2744 508
rect -2944 232 -2744 270
rect -2944 198 -2928 232
rect -2760 198 -2744 232
rect -2944 182 -2744 198
rect -344 522 -144 538
rect -344 488 -328 522
rect -160 488 -144 522
rect -344 450 -144 488
rect -344 212 -144 250
rect -344 178 -328 212
rect -160 178 -144 212
rect -344 162 -144 178
rect 556 742 756 758
rect 556 708 572 742
rect 740 708 756 742
rect 556 670 756 708
rect 556 432 756 470
rect 556 398 572 432
rect 740 398 756 432
rect 556 382 756 398
rect 7796 742 7996 758
rect 7796 708 7812 742
rect 7980 708 7996 742
rect 7796 670 7996 708
rect 7796 432 7996 470
rect 7796 398 7812 432
rect 7980 398 7996 432
rect 7796 382 7996 398
<< polycont >>
rect -5488 3586 -5320 3620
rect -5488 2258 -5320 2292
rect -2928 3586 -2760 3620
rect -2928 2258 -2760 2292
rect -328 3566 -160 3600
rect -328 2238 -160 2272
rect 5932 3346 6100 3380
rect 5932 3018 6100 3052
rect 5932 2426 6100 2460
rect 5932 2098 6100 2132
rect -5488 1646 -5320 1680
rect -5488 918 -5320 952
rect -2928 1626 -2760 1660
rect -2928 898 -2760 932
rect -328 1606 -160 1640
rect -328 878 -160 912
rect 1492 1588 1660 1622
rect 1492 1278 1660 1312
rect 7812 1588 7980 1622
rect 7812 1278 7980 1312
rect -5488 508 -5320 542
rect -5488 198 -5320 232
rect -2928 508 -2760 542
rect -2928 198 -2760 232
rect -328 488 -160 522
rect -328 178 -160 212
rect 572 708 740 742
rect 572 398 740 432
rect 7812 708 7980 742
rect 7812 398 7980 432
<< locali >>
rect -5664 3688 -5568 3722
rect -5240 3688 -5144 3722
rect -5664 3626 -5630 3688
rect -5178 3626 -5144 3688
rect -5504 3586 -5488 3620
rect -5320 3586 -5304 3620
rect -5550 3527 -5516 3543
rect -5550 2335 -5516 2351
rect -5292 3527 -5258 3543
rect -5292 2335 -5258 2351
rect -5504 2258 -5488 2292
rect -5320 2258 -5304 2292
rect -5664 2190 -5630 2252
rect -5178 2190 -5144 2252
rect -5664 2156 -5568 2190
rect -5240 2156 -5144 2190
rect -3104 3688 -3008 3722
rect -2680 3688 -2584 3722
rect -3104 3626 -3070 3688
rect -2618 3626 -2584 3688
rect -2944 3586 -2928 3620
rect -2760 3586 -2744 3620
rect -2990 3527 -2956 3543
rect -2990 2335 -2956 2351
rect -2732 3527 -2698 3543
rect -2732 2335 -2698 2351
rect -2944 2258 -2928 2292
rect -2760 2258 -2744 2292
rect -3104 2190 -3070 2252
rect -2618 2190 -2584 2252
rect -3104 2156 -3008 2190
rect -2680 2156 -2584 2190
rect -504 3668 -408 3702
rect -80 3668 16 3702
rect -504 3606 -470 3668
rect -18 3606 16 3668
rect -344 3566 -328 3600
rect -160 3566 -144 3600
rect -390 3507 -356 3523
rect -390 2315 -356 2331
rect -132 3507 -98 3523
rect -132 2315 -98 2331
rect -344 2238 -328 2272
rect -160 2238 -144 2272
rect -504 2170 -470 2232
rect 5756 3448 5852 3482
rect 6180 3448 6276 3482
rect 5756 3386 5790 3448
rect 6242 3386 6276 3448
rect 5916 3346 5932 3380
rect 6100 3346 6116 3380
rect 5870 3287 5904 3303
rect 5870 3095 5904 3111
rect 6128 3287 6162 3303
rect 6128 3095 6162 3111
rect 5916 3018 5932 3052
rect 6100 3018 6116 3052
rect 5756 2950 5790 3012
rect 6242 2950 6276 3012
rect 5756 2916 5852 2950
rect 6180 2916 6276 2950
rect -18 2170 16 2232
rect -504 2136 -408 2170
rect -80 2136 16 2170
rect 5756 2528 5852 2562
rect 6180 2528 6276 2562
rect 5756 2466 5790 2528
rect 6242 2466 6276 2528
rect 5916 2426 5932 2460
rect 6100 2426 6116 2460
rect 5870 2367 5904 2383
rect 5870 2175 5904 2191
rect 6128 2367 6162 2383
rect 6128 2175 6162 2191
rect 5916 2098 5932 2132
rect 6100 2098 6116 2132
rect 5756 2030 5790 2092
rect 6242 2030 6276 2092
rect 5756 1996 5852 2030
rect 6180 1996 6276 2030
rect -5664 1748 -5568 1782
rect -5240 1748 -5144 1782
rect -5664 1686 -5630 1748
rect -5178 1686 -5144 1748
rect -5504 1646 -5488 1680
rect -5320 1646 -5304 1680
rect -5550 1587 -5516 1603
rect -5550 995 -5516 1011
rect -5292 1587 -5258 1603
rect -5292 995 -5258 1011
rect -5504 918 -5488 952
rect -5320 918 -5304 952
rect -5664 850 -5630 912
rect -5178 850 -5144 912
rect -5664 816 -5568 850
rect -5240 816 -5144 850
rect -3104 1728 -3008 1762
rect -2680 1728 -2584 1762
rect -3104 1666 -3070 1728
rect -2618 1666 -2584 1728
rect -2944 1626 -2928 1660
rect -2760 1626 -2744 1660
rect -2990 1567 -2956 1583
rect -2990 975 -2956 991
rect -2732 1567 -2698 1583
rect -2732 975 -2698 991
rect -2944 898 -2928 932
rect -2760 898 -2744 932
rect -3104 830 -3070 892
rect -2618 830 -2584 892
rect -3104 796 -3008 830
rect -2680 796 -2584 830
rect -504 1708 -408 1742
rect -80 1708 16 1742
rect -504 1646 -470 1708
rect -18 1646 16 1708
rect -344 1606 -328 1640
rect -160 1606 -144 1640
rect -390 1547 -356 1563
rect -390 955 -356 971
rect -132 1547 -98 1563
rect -132 955 -98 971
rect -344 878 -328 912
rect -160 878 -144 912
rect -504 810 -470 872
rect 1316 1690 1412 1724
rect 1740 1690 1836 1724
rect 1316 1628 1350 1690
rect 1802 1628 1836 1690
rect 1476 1588 1492 1622
rect 1660 1588 1676 1622
rect 1430 1538 1464 1554
rect 1430 1346 1464 1362
rect 1688 1538 1722 1554
rect 1688 1346 1722 1362
rect 1476 1278 1492 1312
rect 1660 1278 1676 1312
rect 1316 1210 1350 1272
rect 1802 1210 1836 1272
rect 1316 1176 1412 1210
rect 1740 1176 1836 1210
rect 7636 1690 7732 1724
rect 8060 1690 8156 1724
rect 7636 1628 7670 1690
rect 8122 1628 8156 1690
rect 7796 1588 7812 1622
rect 7980 1588 7996 1622
rect 7750 1538 7784 1554
rect 7750 1346 7784 1362
rect 8008 1538 8042 1554
rect 8008 1346 8042 1362
rect 7796 1278 7812 1312
rect 7980 1278 7996 1312
rect 7636 1210 7670 1272
rect 8122 1210 8156 1272
rect 7636 1176 7732 1210
rect 8060 1176 8156 1210
rect -18 810 16 872
rect -504 776 -408 810
rect -80 776 16 810
rect 396 810 492 844
rect 820 810 916 844
rect 396 748 430 810
rect -5664 610 -5568 644
rect -5240 610 -5144 644
rect -5664 548 -5630 610
rect -5178 548 -5144 610
rect -5504 508 -5488 542
rect -5320 508 -5304 542
rect -5550 458 -5516 474
rect -5550 266 -5516 282
rect -5292 458 -5258 474
rect -5292 266 -5258 282
rect -5504 198 -5488 232
rect -5320 198 -5304 232
rect -5664 130 -5630 192
rect -5178 130 -5144 192
rect -5664 96 -5568 130
rect -5240 96 -5144 130
rect -3104 610 -3008 644
rect -2680 610 -2584 644
rect -3104 548 -3070 610
rect -2618 548 -2584 610
rect -2944 508 -2928 542
rect -2760 508 -2744 542
rect -2990 458 -2956 474
rect -2990 266 -2956 282
rect -2732 458 -2698 474
rect -2732 266 -2698 282
rect -2944 198 -2928 232
rect -2760 198 -2744 232
rect -3104 130 -3070 192
rect -2618 130 -2584 192
rect -3104 96 -3008 130
rect -2680 96 -2584 130
rect -504 590 -408 624
rect -80 590 16 624
rect -504 528 -470 590
rect -18 528 16 590
rect -344 488 -328 522
rect -160 488 -144 522
rect -390 438 -356 454
rect -390 246 -356 262
rect -132 438 -98 454
rect -132 246 -98 262
rect -344 178 -328 212
rect -160 178 -144 212
rect -504 110 -470 172
rect 882 748 916 810
rect 556 708 572 742
rect 740 708 756 742
rect 510 658 544 674
rect 510 466 544 482
rect 768 658 802 674
rect 768 466 802 482
rect 556 398 572 432
rect 740 398 756 432
rect 396 330 430 392
rect 882 330 916 392
rect 396 296 492 330
rect 820 296 916 330
rect 7636 810 7732 844
rect 8060 810 8156 844
rect 7636 748 7670 810
rect 8122 748 8156 810
rect 7796 708 7812 742
rect 7980 708 7996 742
rect 7750 658 7784 674
rect 7750 466 7784 482
rect 8008 658 8042 674
rect 8008 466 8042 482
rect 7796 398 7812 432
rect 7980 398 7996 432
rect 7636 330 7670 392
rect 8122 330 8156 392
rect 7636 296 7732 330
rect 8060 296 8156 330
rect -18 110 16 172
rect -504 76 -408 110
rect -80 76 16 110
<< metal1 >>
rect -1660 4154 -1550 4250
rect -3811 3954 149 4154
rect -1210 3570 -150 3710
rect -6380 2380 -5025 2490
rect -290 2200 -150 3570
rect -51 2687 149 3954
rect -290 2100 -280 2200
rect -160 2100 -150 2200
rect -290 2090 -150 2100
rect -6380 1660 -5130 1800
rect -613 1694 136 1894
rect -300 1500 -140 1520
rect -300 1400 -280 1500
rect -160 1400 -140 1500
rect -300 980 -140 1400
rect -6380 760 -5220 920
rect -300 820 100 980
rect 8120 780 8260 920
rect 1840 20 2220 40
rect -6420 -60 -5300 -40
rect -6420 -220 -6160 -60
rect -6020 -220 -5300 -60
rect -6420 -240 -5300 -220
rect 1840 -220 1860 20
rect 2200 -220 2220 20
rect 1840 -240 2220 -220
<< via1 >>
rect -280 2100 -160 2200
rect -280 1400 -160 1500
rect -6160 -220 -6020 -60
rect 1860 -220 2200 20
<< metal2 >>
rect -300 2200 -140 2220
rect -300 2100 -280 2200
rect -160 2100 -140 2200
rect -300 2080 -140 2100
rect -280 1520 -160 2080
rect -300 1500 -140 1520
rect -300 1400 -280 1500
rect -160 1400 -140 1500
rect -300 1380 -140 1400
rect -2780 390 -2600 400
rect -2780 210 810 390
rect -2780 -40 -2600 210
rect 630 -40 810 210
rect 1840 20 2220 40
rect 1840 -40 1860 20
rect -6180 -60 -5940 -40
rect -6180 -220 -6160 -60
rect -6020 -220 -5940 -60
rect -6180 -240 -5940 -220
rect -4940 -240 -2000 -40
rect 620 -220 1860 -40
rect 2200 -220 2220 20
rect 620 -240 2220 -220
use buffer  buffer_0 ~/projects-sky130/temp-sensor/amp-op/mag/buffer
timestamp 1668731387
transform 1 0 -13880 0 1 -1424
box 13875 1430 22120 4938
use ota  ota_0 ~/projects-sky130/temp-sensor/amp-op/mag/ota
timestamp 1668746219
transform 1 0 -4851 0 1 -4906
box -540 140 4440 9060
<< labels >>
flabel metal1 -6380 760 -6220 920 0 FreeSans 1600 0 0 0 in2
port 9 nsew
flabel metal1 -6400 -240 -6200 -60 0 FreeSans 1600 0 0 0 vs
port 5 nsew
flabel metal1 -6380 1660 -6220 1800 0 FreeSans 1600 0 0 0 in1
port 3 nsew
flabel metal1 -6380 2380 -6270 2490 0 FreeSans 1600 0 0 0 ib
port 2 nsew
flabel metal1 8120 780 8260 920 0 FreeSans 1600 0 0 0 out
port 7 nsew
flabel metal1 -1660 4140 -1550 4250 0 FreeSans 1600 0 0 0 vd
port 1 nsew
<< end >>
