** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex_tb-ac.sch
**.subckt impedance-transformer-pex_tb-ac
Vin net1 GND DC 0 AC 1
Vin1 net2 GND DC 0 AC 1
R3 ns12 GND 50 m=1
R4 ns22 net2 50 m=1
xit1 ns11 ns12 GND impedance-transformer-pex
xit2 ns21 ns22 GND impedance-transformer-pex
R1 net1 ns11 172.7 m=1
R2 GND ns21 172.7 m=1
**** begin user architecture code



.ac lin 1MEG 1.5G 4G
.control
destroy all
set units=degrees
run

set color0=white
set color1=black

let z0=50
let zl=169

* Find two S parameters from test circuit
let s11 = v(ns11)
let s12 = v(ns12)
let s21 = v(ns21)
let s22 = v(ns22)

* Extract Y parameters
*let StoYDelS = ((1+s11)*(1+s22)-s12*s21)*z0
*let y11 = ((1+s22)*(1-s11)+s12*s21/StoYDelS
*let y12=-2*s12/StoYDelS
*let y21=-2*s21/StoYDelS
*let y22 = ((1+s11)*(1-s22)+s12+s21)/StoYDelS

* Extract Z parameters
let StoZDelS = ((1-s11)*(1-s22)-s12*s21)/z0
let z11 = ((1+s11)*(1-s22)+s12*s21)/StoZDelS
let z12 = 2*s12/StoZDelS
let z21 = 2*s21/StoZDelS
let z22=((1-s11)*(1+s22)+s12*s21)/StoZDelS

*plot z11
*plot z12
*plot z21
*plot z22 xlimit 2.4G 2.5G
*plot ph(z22) xlimit 2.4G 2.5G
*plot z22
*plot smith z22
let z_in =z11-z12*z21/(z22+z0)
plot ph(z_in)
plot mag(z_in)
let z_output=z22-(z12*z21/(z11+zl))
plot ph(z_output)
plot mag(z_output)
let gamma=(mag(z_output)-mag(z_in))/(mag(z_output)+mag(z_in))
plot gamma*100
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex.sym # of pins=3
** sym_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex.sym
** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex.sch
.subckt impedance-transformer-pex  in out gnd
*.iopin gnd
*.iopin in
*.iopin out
xl1 in out l1
**** begin user architecture code

* NGSPICE file created from impedance-transformer.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_2_3YFQRG m4_n2675_n10534# c2_n2575_n10434# VSUBS
X0 c2_n2575_n10434# m4_n2675_n10534# sky130_fd_pr__cap_mim_m3_2 l=2.496e+07u w=2.496e+07u
X1 c2_n2575_n10434# m4_n2675_n10534# sky130_fd_pr__cap_mim_m3_2 l=2.496e+07u w=2.496e+07u
X2 c2_n2575_n10434# m4_n2675_n10534# sky130_fd_pr__cap_mim_m3_2 l=2.496e+07u w=2.496e+07u
X3 c2_n2575_n10434# m4_n2675_n10534# sky130_fd_pr__cap_mim_m3_2 l=2.496e+07u w=2.496e+07u
C0 c2_n2575_n10434# m4_n2675_n10534# 164.66fF
C1 c2_n2575_n10434# VSUBS 0.30fF
C2 m4_n2675_n10534# VSUBS 42.24fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_93FFAE c2_n2522_n7629# m4_n2622_n7729# VSUBS
X0 c2_n2522_n7629# m4_n2622_n7729# sky130_fd_pr__cap_mim_m3_2 l=2.443e+07u w=2.443e+07u
X1 c2_n2522_n7629# m4_n2622_n7729# sky130_fd_pr__cap_mim_m3_2 l=2.443e+07u w=2.443e+07u
X2 c2_n2522_n7629# m4_n2622_n7729# sky130_fd_pr__cap_mim_m3_2 l=2.443e+07u w=2.443e+07u
C0 c2_n2522_n7629# m4_n2622_n7729# 118.74fF
C1 c2_n2522_n7629# VSUBS 0.26fF
C2 m4_n2622_n7729# VSUBS 30.75fF
.ends

*.subckt impedance-transformer gnd out in
Xsky130_fd_pr__cap_mim_m3_2_3YFQRG_0 gnd out gnd sky130_fd_pr__cap_mim_m3_2_3YFQRG
Xsky130_fd_pr__cap_mim_m3_2_3YFQRG_1 gnd out gnd sky130_fd_pr__cap_mim_m3_2_3YFQRG
Xsky130_fd_pr__cap_mim_m3_2_3YFQRG_2 gnd out gnd sky130_fd_pr__cap_mim_m3_2_3YFQRG
Xsky130_fd_pr__cap_mim_m3_2_3YFQRG_3 gnd out gnd sky130_fd_pr__cap_mim_m3_2_3YFQRG
Xsky130_fd_pr__cap_mim_m3_2_93FFAE_0 in gnd gnd sky130_fd_pr__cap_mim_m3_2_93FFAE
Xsky130_fd_pr__cap_mim_m3_2_93FFAE_1 in gnd gnd sky130_fd_pr__cap_mim_m3_2_93FFAE
Xsky130_fd_pr__cap_mim_m3_2_93FFAE_2 in gnd gnd sky130_fd_pr__cap_mim_m3_2_93FFAE

R0 out out.n2 0.192
R1 out.t15 out.t13 0.066
R2 out.t14 out.t15 0.066
R3 out.t12 out.t14 0.066
R4 out.t11 out.t9 0.066
R5 out.t10 out.t11 0.066
R6 out.t8 out.t10 0.066
R7 out.t7 out.t5 0.066
R8 out.t6 out.t7 0.066
R9 out.t4 out.t6 0.066
R10 out.t3 out.t1 0.066
R11 out.t2 out.t3 0.066
R12 out.t0 out.t2 0.066
R13 out.n1 out.t0 0.062
R14 out.n0 out.t12 0.056
R15 out.n1 out.t4 0.047
R16 out.n0 out.t8 0.046
R17 out.n2 out.n1 0.006
R18 out.n2 out.n0 0.004
R19 in in.n0 0.26
R20 in.t2 in.t0 0.066
R21 in.t1 in.t2 0.066
R22 in.t5 in.t3 0.066
R23 in.t4 in.t5 0.066
R24 in.t8 in.t6 0.066
R25 in.t7 in.t8 0.064
R26 in.n0 in.t1 0.05
R27 in.n0 in.t7 0.047
R28 in.n0 in.t4 0.039
C0 in.t6 gnd 14.51fF
C1 in.t8 gnd 14.50fF
C2 in.t7 gnd 37.65fF
C3 in.t3 gnd 14.51fF
C4 in.t5 gnd 14.54fF
C5 in.t4 gnd 14.38fF
C6 in.t0 gnd 14.51fF
C7 in.t2 gnd 14.54fF
C8 in.t1 gnd 20.60fF
C9 in.n0 gnd 474.44fF $ **FLOATING
C10 out.t9 gnd 17.89fF
C11 out.t11 gnd 17.93fF
C12 out.t10 gnd 17.93fF
C13 out.t8 gnd 18.23fF
C14 out.t13 gnd 17.89fF
C15 out.t15 gnd 17.93fF
C16 out.t14 gnd 17.93fF
C17 out.t12 gnd 24.02fF
C18 out.n0 gnd 54.72fF $ **FLOATING
C19 out.t5 gnd 17.89fF
C20 out.t7 gnd 17.93fF
C21 out.t6 gnd 17.93fF
C22 out.t4 gnd 18.28fF
C23 out.t1 gnd 17.89fF
C24 out.t3 gnd 17.93fF
C25 out.t2 gnd 17.93fF
C26 out.t0 gnd 22.51fF
C27 out.n1 gnd 54.23fF $ **FLOATING
C28 out.n2 gnd 512.64fF $ **FLOATING
C29 in gnd 311.92fF
C30 out gnd 306.12fF
*.ends



**** end user architecture code
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sym
*+ # of pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sch
.subckt l1  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 592.7p m=1
Cs1 p1 net1 26.83f m=1
Cs2 p2 net2 24.25f m=1
Rs1 net1 GND 65.02 m=1
Rs2 net2 GND 14.4 m=1
R1 p2 net3 2.935 m=1
.ends

.GLOBAL GND
.end
