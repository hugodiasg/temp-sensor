magic
tech sky130A
magscale 1 2
timestamp 1647142466
<< error_p >>
rect -2586 5164 2586 5304
rect -2586 4924 2586 5064
rect -2586 50 2586 190
rect -2586 -190 2586 -50
rect -2586 -5064 2586 -4924
rect -2586 -5304 2586 -5164
<< metal4 >>
rect -2586 10137 2586 10178
rect -2586 5205 2330 10137
rect 2566 5205 2586 10137
rect -2586 5164 2586 5205
rect -2586 5023 2586 5064
rect -2586 91 2330 5023
rect 2566 91 2586 5023
rect -2586 50 2586 91
rect -2586 -91 2586 -50
rect -2586 -5023 2330 -91
rect 2566 -5023 2586 -91
rect -2586 -5064 2586 -5023
rect -2586 -5205 2586 -5164
rect -2586 -10137 2330 -5205
rect 2566 -10137 2586 -5205
rect -2586 -10178 2586 -10137
<< via4 >>
rect 2330 5205 2566 10137
rect 2330 91 2566 5023
rect 2330 -5023 2566 -91
rect 2330 -10137 2566 -5205
<< mimcap2 >>
rect -2486 10038 2328 10078
rect -2486 5304 -1973 10038
rect 1815 5304 2328 10038
rect -2486 5264 2328 5304
rect -2486 4924 2328 4964
rect -2486 190 -1973 4924
rect 1815 190 2328 4924
rect -2486 150 2328 190
rect -2486 -190 2328 -150
rect -2486 -4924 -1973 -190
rect 1815 -4924 2328 -190
rect -2486 -4964 2328 -4924
rect -2486 -5304 2328 -5264
rect -2486 -10038 -1973 -5304
rect 1815 -10038 2328 -5304
rect -2486 -10078 2328 -10038
<< mimcap2contact >>
rect -1973 5304 1815 10038
rect -1973 190 1815 4924
rect -1973 -4924 1815 -190
rect -1973 -10038 1815 -5304
<< metal5 >>
rect -239 10062 81 10228
rect 2288 10137 2608 10228
rect -1997 10038 1839 10062
rect -1997 5304 -1973 10038
rect 1815 5304 1839 10038
rect -1997 5280 1839 5304
rect -239 4948 81 5280
rect 2288 5205 2330 10137
rect 2566 5205 2608 10137
rect 2288 5023 2608 5205
rect -1997 4924 1839 4948
rect -1997 190 -1973 4924
rect 1815 190 1839 4924
rect -1997 166 1839 190
rect -239 -166 81 166
rect 2288 91 2330 5023
rect 2566 91 2608 5023
rect 2288 -91 2608 91
rect -1997 -190 1839 -166
rect -1997 -4924 -1973 -190
rect 1815 -4924 1839 -190
rect -1997 -4948 1839 -4924
rect -239 -5280 81 -4948
rect 2288 -5023 2330 -91
rect 2566 -5023 2608 -91
rect 2288 -5205 2608 -5023
rect -1997 -5304 1839 -5280
rect -1997 -10038 -1973 -5304
rect 1815 -10038 1839 -5304
rect -1997 -10062 1839 -10038
rect -239 -10228 81 -10062
rect 2288 -10137 2330 -5205
rect 2566 -10137 2608 -5205
rect 2288 -10228 2608 -10137
<< properties >>
string FIXED_BBOX -2586 5164 2428 10178
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.07 l 24.07 val 1.177k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
