magic
tech sky130A
magscale 1 2
timestamp 1643981260
<< metal4 >>
rect -2801 2509 2801 2550
rect -2801 -2509 2545 2509
rect 2781 -2509 2801 2509
rect -2801 -2550 2801 -2509
<< via4 >>
rect 2545 -2509 2781 2509
<< mimcap2 >>
rect -2701 2410 2199 2450
rect -2701 -2410 -2661 2410
rect 2159 -2410 2199 2410
rect -2701 -2450 2199 -2410
<< mimcap2contact >>
rect -2661 -2410 2159 2410
<< metal5 >>
rect 2503 2509 2823 2551
rect -2685 2410 2183 2434
rect -2685 -2410 -2661 2410
rect 2159 -2410 2183 2410
rect -2685 -2434 2183 -2410
rect 2503 -2509 2545 2509
rect 2781 -2509 2823 2509
rect 2503 -2551 2823 -2509
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2801 -2550 2299 2550
string parameters w 24.5 l 24.5 val 1.219k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
