magic
tech sky130
timestamp 1643667960
<< checkpaint >>
rect -2125 -2075 2124 2075
<< metal3 >>
rect -2125 -2075 2124 -2047
rect -2125 -2047 2040 2047
rect 2104 -2047 2124 2047
rect -2125 2047 2124 2075
<< via3 >>
rect 2040 -2047 2104 2047
<< metal4 >>
rect -1986 -1936 1886 -1935
rect -1986 -1935 -1985 1935
rect 1885 -1935 1886 1935
rect -1986 1935 1886 1936
rect 2024 -2063 2120 -2047
rect 2024 -2047 2040 2047
rect 2104 -2047 2120 2047
rect 2024 2047 2120 2063
<< mimcap >>
rect -2025 -1975 1925 -1935
rect -2025 -1935 -1985 1935
rect 1885 -1935 1925 1935
rect -2025 1935 1925 1975
<< mimcapcontact >>
rect -1985 -1935 1885 1935
<< end >>
