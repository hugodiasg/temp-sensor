magic
tech sky130A
magscale 1 2
timestamp 1668746219
<< psubdiff >>
rect -424 4400 -400 4540
rect -200 4400 -176 4540
<< psubdiffcont >>
rect -400 4400 -200 4540
<< viali >>
rect -420 4400 -400 4540
rect -400 4400 -200 4540
rect -200 4400 -180 4540
<< metal1 >>
rect 1040 8860 1240 9060
rect 600 8700 1620 8860
rect 200 8600 340 8620
rect 200 8500 220 8600
rect 320 8500 340 8600
rect 200 8480 340 8500
rect 600 8440 760 8700
rect 1060 8600 1200 8620
rect 1060 8500 1080 8600
rect 1180 8500 1200 8600
rect 1060 8480 1200 8500
rect 400 8280 760 8440
rect 1460 8420 1620 8700
rect 2860 8600 3000 8620
rect 2860 8500 2880 8600
rect 2980 8500 3000 8600
rect 2860 8480 3000 8500
rect 3140 8600 3280 8620
rect 3140 8500 3160 8600
rect 3260 8500 3280 8600
rect 3140 8480 3280 8500
rect 3400 8600 3540 8620
rect 3400 8500 3420 8600
rect 3520 8500 3540 8600
rect 3400 8480 3540 8500
rect 3640 8600 3780 8620
rect 3640 8500 3660 8600
rect 3760 8500 3780 8600
rect 3640 8480 3780 8500
rect 1280 8280 3880 8420
rect 3040 7560 3620 7580
rect -540 7260 340 7460
rect 40 7160 340 7260
rect 640 7260 1040 7460
rect 3040 7360 4240 7560
rect -540 6540 380 6740
rect 640 6500 840 7260
rect 4040 6800 4240 7360
rect 4040 6600 4440 6800
rect -540 5820 -140 5840
rect -540 5660 -320 5820
rect -160 5660 -140 5820
rect -540 5640 -140 5660
rect -20 5560 160 6480
rect 420 6300 1040 6500
rect 1300 6340 3580 6540
rect 1020 5820 1220 5840
rect 1020 5660 1040 5820
rect 1200 5660 1220 5820
rect 1020 5640 1220 5660
rect -20 5420 1240 5560
rect -20 5200 160 5420
rect 420 5200 1020 5380
rect 1300 5360 1700 6340
rect 4040 6280 4240 6600
rect 3040 6080 4240 6280
rect 1300 5220 1520 5360
rect 1660 5220 1700 5360
rect 1300 5200 1700 5220
rect 2690 5550 3390 5730
rect 2690 5240 2870 5550
rect 630 5050 810 5200
rect 2690 5140 3680 5240
rect 90 4860 1350 5050
rect 2690 4860 2870 5140
rect 4040 5000 4240 6080
rect -540 4670 2870 4860
rect 3380 4980 4240 5000
rect 3380 4820 3400 4980
rect 3620 4820 4240 4980
rect 3380 4800 4240 4820
rect -540 4660 2860 4670
rect -440 4540 -160 4660
rect -440 4400 -420 4540
rect -180 4400 -160 4540
rect -440 4380 -160 4400
<< via1 >>
rect 220 8500 320 8600
rect 1080 8500 1180 8600
rect 2880 8500 2980 8600
rect 3160 8500 3260 8600
rect 3420 8500 3520 8600
rect 3660 8500 3760 8600
rect -320 5660 -160 5820
rect 1040 5660 1200 5820
rect 1520 5220 1660 5360
rect 3400 4820 3620 4980
<< metal2 >>
rect 180 8600 3880 8680
rect 180 8500 220 8600
rect 320 8500 1080 8600
rect 1180 8500 2880 8600
rect 2980 8500 3160 8600
rect 3260 8500 3420 8600
rect 3520 8500 3660 8600
rect 3760 8500 3880 8600
rect 180 8480 3880 8500
rect -340 5820 1220 5840
rect -340 5660 -320 5820
rect -160 5660 1040 5820
rect 1200 5660 1220 5820
rect -340 5640 1220 5660
rect 1500 5360 1680 5380
rect 1500 5220 1520 5360
rect 1660 5220 1680 5360
rect 1500 5200 1680 5220
rect 3380 4980 3640 5000
rect 3380 4820 3400 4980
rect 3620 4820 3640 4980
rect 3380 4800 3640 4820
<< via2 >>
rect 1520 5220 1660 5360
rect 3400 4820 3620 4980
<< metal3 >>
rect 1500 5360 1700 5380
rect 1500 5220 1520 5360
rect 1660 5220 1700 5360
rect 1500 4340 1700 5220
rect 3380 4980 3640 5000
rect 3380 4820 3400 4980
rect 3620 4820 3640 4980
rect 3380 4800 3640 4820
<< via3 >>
rect 3400 4820 3620 4980
<< metal4 >>
rect 3380 4980 3640 5000
rect 3380 4820 3400 4980
rect 3620 4820 3640 4980
rect 3380 4180 3640 4820
use sky130_fd_pr__cap_mim_m3_1_2NYK3R  XCC
timestamp 1668740706
transform 1 0 2170 0 1 2340
box -2250 -2200 2249 2200
use sky130_fd_pr__pfet_01v8_G8TFUZ  XM1
timestamp 1668740706
transform 1 0 296 0 1 6199
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_G8PDUZ  XM2
timestamp 1668741396
transform 1 0 1156 0 1 6199
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_SXTBPF  XM4
timestamp 1668741396
transform 1 0 1157 0 1 5291
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_G8TPYT  XM5
timestamp 1668740706
transform 1 0 296 0 1 7839
box -296 -819 296 819
use sky130_fd_pr__nfet_01v8_XABGW3  XM7
timestamp 1668741396
transform 1 0 3345 0 1 5840
box -425 -660 425 660
use sky130_fd_pr__pfet_01v8_8ALGB7  XM8
timestamp 1668740706
transform 1 0 3343 0 1 7689
box -683 -969 683 969
use sky130_fd_pr__nfet_01v8_SXTBPF  sky130_fd_pr__nfet_01v8_SXTBPF_0
timestamp 1668741396
transform 1 0 297 0 1 5291
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_G8TPYT  sky130_fd_pr__pfet_01v8_G8TPYT_0
timestamp 1668740706
transform 1 0 1156 0 1 7839
box -296 -819 296 819
<< labels >>
flabel metal1 1040 8860 1240 9060 0 FreeSans 128 0 0 0 vd
port 0 nsew
flabel metal1 4240 6600 4440 6800 0 FreeSans 128 0 0 0 out
port 5 nsew
flabel metal1 -540 7260 -340 7460 0 FreeSans 128 0 0 0 ib
port 2 nsew
flabel metal1 -540 6540 -340 6740 0 FreeSans 128 0 0 0 in1
port 3 nsew
flabel metal1 -540 5640 -340 5840 0 FreeSans 128 0 0 0 in2
port 4 nsew
flabel metal1 -540 4660 -340 4860 0 FreeSans 128 0 0 0 vs
port 1 nsew
<< end >>
