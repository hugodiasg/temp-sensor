magic
tech sky130A
magscale 1 2
timestamp 1645495691
<< metal4 >>
rect -2635 7727 2635 7768
rect -2635 2697 2379 7727
rect 2615 2697 2635 7727
rect -2635 2656 2635 2697
rect -2635 2515 2635 2556
rect -2635 -2515 2379 2515
rect 2615 -2515 2635 2515
rect -2635 -2556 2635 -2515
rect -2635 -2697 2635 -2656
rect -2635 -7727 2379 -2697
rect 2615 -7727 2635 -2697
rect -2635 -7768 2635 -7727
<< via4 >>
rect 2379 2697 2615 7727
rect 2379 -2515 2615 2515
rect 2379 -7727 2615 -2697
<< mimcap2 >>
rect -2535 7628 2377 7668
rect -2535 2796 -2012 7628
rect 1854 2796 2377 7628
rect -2535 2756 2377 2796
rect -2535 2416 2377 2456
rect -2535 -2416 -2012 2416
rect 1854 -2416 2377 2416
rect -2535 -2456 2377 -2416
rect -2535 -2796 2377 -2756
rect -2535 -7628 -2012 -2796
rect 1854 -7628 2377 -2796
rect -2535 -7668 2377 -7628
<< mimcap2contact >>
rect -2012 2796 1854 7628
rect -2012 -2416 1854 2416
rect -2012 -7628 1854 -2796
<< metal5 >>
rect -239 7652 81 7818
rect 2337 7727 2657 7818
rect -2036 7628 1878 7652
rect -2036 2796 -2012 7628
rect 1854 2796 1878 7628
rect -2036 2772 1878 2796
rect -239 2440 81 2772
rect 2337 2697 2379 7727
rect 2615 2697 2657 7727
rect 2337 2515 2657 2697
rect -2036 2416 1878 2440
rect -2036 -2416 -2012 2416
rect 1854 -2416 1878 2416
rect -2036 -2440 1878 -2416
rect -239 -2772 81 -2440
rect 2337 -2515 2379 2515
rect 2615 -2515 2657 2515
rect 2337 -2697 2657 -2515
rect -2036 -2796 1878 -2772
rect -2036 -7628 -2012 -2796
rect 1854 -7628 1878 -2796
rect -2036 -7652 1878 -7628
rect -239 -7818 81 -7652
rect 2337 -7727 2379 -2697
rect 2615 -7727 2657 -2697
rect 2337 -7818 2657 -7727
<< properties >>
string FIXED_BBOX -2635 2656 2477 7768
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.559 l 24.559 val 1.224k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
