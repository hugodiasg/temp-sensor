magic
tech sky130A
timestamp 1643669011
<< pwell >>
rect -422 -339 422 339
<< mvnmos >>
rect -308 -210 -208 210
rect -179 -210 -79 210
rect -50 -210 50 210
rect 79 -210 179 210
rect 208 -210 308 210
<< mvndiff >>
rect -337 204 -308 210
rect -337 -204 -331 204
rect -314 -204 -308 204
rect -337 -210 -308 -204
rect -208 204 -179 210
rect -208 -204 -202 204
rect -185 -204 -179 204
rect -208 -210 -179 -204
rect -79 204 -50 210
rect -79 -204 -73 204
rect -56 -204 -50 204
rect -79 -210 -50 -204
rect 50 204 79 210
rect 50 -204 56 204
rect 73 -204 79 204
rect 50 -210 79 -204
rect 179 204 208 210
rect 179 -204 185 204
rect 202 -204 208 204
rect 179 -210 208 -204
rect 308 204 337 210
rect 308 -204 314 204
rect 331 -204 337 204
rect 308 -210 337 -204
<< mvndiffc >>
rect -331 -204 -314 204
rect -202 -204 -185 204
rect -73 -204 -56 204
rect 56 -204 73 204
rect 185 -204 202 204
rect 314 -204 331 204
<< mvpsubdiff >>
rect -404 315 404 321
rect -404 298 -350 315
rect 350 298 404 315
rect -404 292 404 298
rect -404 267 -375 292
rect -404 -267 -398 267
rect -381 -267 -375 267
rect 375 267 404 292
rect -404 -292 -375 -267
rect 375 -267 381 267
rect 398 -267 404 267
rect 375 -292 404 -267
rect -404 -298 404 -292
rect -404 -315 -350 -298
rect 350 -315 404 -298
rect -404 -321 404 -315
<< mvpsubdiffcont >>
rect -350 298 350 315
rect -398 -267 -381 267
rect 381 -267 398 267
rect -350 -315 350 -298
<< poly >>
rect -308 246 -208 254
rect -308 229 -300 246
rect -216 229 -208 246
rect -308 210 -208 229
rect -179 246 -79 254
rect -179 229 -171 246
rect -87 229 -79 246
rect -179 210 -79 229
rect -50 246 50 254
rect -50 229 -42 246
rect 42 229 50 246
rect -50 210 50 229
rect 79 246 179 254
rect 79 229 87 246
rect 171 229 179 246
rect 79 210 179 229
rect 208 246 308 254
rect 208 229 216 246
rect 300 229 308 246
rect 208 210 308 229
rect -308 -229 -208 -210
rect -308 -246 -300 -229
rect -216 -246 -208 -229
rect -308 -254 -208 -246
rect -179 -229 -79 -210
rect -179 -246 -171 -229
rect -87 -246 -79 -229
rect -179 -254 -79 -246
rect -50 -229 50 -210
rect -50 -246 -42 -229
rect 42 -246 50 -229
rect -50 -254 50 -246
rect 79 -229 179 -210
rect 79 -246 87 -229
rect 171 -246 179 -229
rect 79 -254 179 -246
rect 208 -229 308 -210
rect 208 -246 216 -229
rect 300 -246 308 -229
rect 208 -254 308 -246
<< polycont >>
rect -300 229 -216 246
rect -171 229 -87 246
rect -42 229 42 246
rect 87 229 171 246
rect 216 229 300 246
rect -300 -246 -216 -229
rect -171 -246 -87 -229
rect -42 -246 42 -229
rect 87 -246 171 -229
rect 216 -246 300 -229
<< locali >>
rect -398 298 -350 315
rect 350 298 398 315
rect -398 267 -381 298
rect 381 267 398 298
rect -308 229 -300 246
rect -216 229 -208 246
rect -179 229 -171 246
rect -87 229 -79 246
rect -50 229 -42 246
rect 42 229 50 246
rect 79 229 87 246
rect 171 229 179 246
rect 208 229 216 246
rect 300 229 308 246
rect -331 204 -314 212
rect -331 -212 -314 -204
rect -202 204 -185 212
rect -202 -212 -185 -204
rect -73 204 -56 212
rect -73 -212 -56 -204
rect 56 204 73 212
rect 56 -212 73 -204
rect 185 204 202 212
rect 185 -212 202 -204
rect 314 204 331 212
rect 314 -212 331 -204
rect -308 -246 -300 -229
rect -216 -246 -208 -229
rect -179 -246 -171 -229
rect -87 -246 -79 -229
rect -50 -246 -42 -229
rect 42 -246 50 -229
rect 79 -246 87 -229
rect 171 -246 179 -229
rect 208 -246 216 -229
rect 300 -246 308 -229
rect -398 -315 -381 -267
rect 381 -315 398 -267
<< viali >>
rect -300 229 -216 246
rect -171 229 -87 246
rect -42 229 42 246
rect 87 229 171 246
rect 216 229 300 246
rect -331 -204 -314 204
rect -202 -204 -185 204
rect -73 -204 -56 204
rect 56 -204 73 204
rect 185 -204 202 204
rect 314 -204 331 204
rect -300 -246 -216 -229
rect -171 -246 -87 -229
rect -42 -246 42 -229
rect 87 -246 171 -229
rect 216 -246 300 -229
rect -381 -315 -350 -298
rect -350 -315 350 -298
rect 350 -315 381 -298
<< metal1 >>
rect -306 246 -210 249
rect -306 229 -300 246
rect -216 229 -210 246
rect -306 226 -210 229
rect -177 246 -81 249
rect -177 229 -171 246
rect -87 229 -81 246
rect -177 226 -81 229
rect -48 246 48 249
rect -48 229 -42 246
rect 42 229 48 246
rect -48 226 48 229
rect 81 246 177 249
rect 81 229 87 246
rect 171 229 177 246
rect 81 226 177 229
rect 210 246 306 249
rect 210 229 216 246
rect 300 229 306 246
rect 210 226 306 229
rect -334 204 -311 210
rect -334 -204 -331 204
rect -314 -204 -311 204
rect -334 -210 -311 -204
rect -205 204 -182 210
rect -205 -204 -202 204
rect -185 -204 -182 204
rect -205 -210 -182 -204
rect -76 204 -53 210
rect -76 -204 -73 204
rect -56 -204 -53 204
rect -76 -210 -53 -204
rect 53 204 76 210
rect 53 -204 56 204
rect 73 -204 76 204
rect 53 -210 76 -204
rect 182 204 205 210
rect 182 -204 185 204
rect 202 -204 205 204
rect 182 -210 205 -204
rect 311 204 334 210
rect 311 -204 314 204
rect 331 -204 334 204
rect 311 -210 334 -204
rect -306 -229 -210 -226
rect -306 -246 -300 -229
rect -216 -246 -210 -229
rect -306 -249 -210 -246
rect -177 -229 -81 -226
rect -177 -246 -171 -229
rect -87 -246 -81 -229
rect -177 -249 -81 -246
rect -48 -229 48 -226
rect -48 -246 -42 -229
rect 42 -246 48 -229
rect -48 -249 48 -246
rect 81 -229 177 -226
rect 81 -246 87 -229
rect 171 -246 177 -229
rect 81 -249 177 -246
rect 210 -229 306 -226
rect 210 -246 216 -229
rect 300 -246 306 -229
rect 210 -249 306 -246
rect -387 -298 387 -295
rect -387 -315 -381 -298
rect 381 -315 387 -298
rect -387 -318 387 -315
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -389 -306 389 306
string parameters w 4.2 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
