magic
tech sky130A
magscale 1 2
timestamp 1644161670
<< error_p >>
rect 1942 2716 1979 7484
rect 1942 -2384 1979 2384
rect 1942 -7484 1979 -2716
rect 2262 -7650 2299 7650
rect 2582 2599 2619 2821
rect 2582 2279 2619 2501
rect 2582 -2501 2619 -2279
rect 2582 -2821 2619 -2599
<< metal4 >>
rect -2598 7559 2597 7600
rect -2598 2641 2341 7559
rect 2577 2641 2597 7559
rect -2598 2600 2597 2641
rect -2598 2459 2597 2500
rect -2598 -2459 2341 2459
rect 2577 -2459 2597 2459
rect -2598 -2500 2597 -2459
rect -2598 -2641 2597 -2600
rect -2598 -7559 2341 -2641
rect 2577 -7559 2597 -2641
rect -2598 -7600 2597 -7559
<< via4 >>
rect 2341 2641 2577 7559
rect 2341 -2459 2577 2459
rect 2341 -7559 2577 -2641
<< mimcap2 >>
rect -2498 7460 2302 7500
rect -2498 2740 -2151 7460
rect 1955 2740 2302 7460
rect -2498 2700 2302 2740
rect -2498 2360 2302 2400
rect -2498 -2360 -2151 2360
rect 1955 -2360 2302 2360
rect -2498 -2400 2302 -2360
rect -2498 -2740 2302 -2700
rect -2498 -7460 -2151 -2740
rect 1955 -7460 2302 -2740
rect -2498 -7500 2302 -7460
<< mimcap2contact >>
rect -2151 2740 1955 7460
rect -2151 -2360 1955 2360
rect -2151 -7460 1955 -2740
<< metal5 >>
rect -258 7484 62 7650
rect 2262 7601 2582 7650
rect 2262 7559 2619 7601
rect -2175 7460 1979 7484
rect -2175 2740 -2151 7460
rect 1955 2740 1979 7460
rect -2175 2716 1979 2740
rect -258 2384 62 2716
rect 2262 2641 2341 7559
rect 2577 2641 2619 7559
rect 2262 2599 2619 2641
rect 2262 2501 2582 2599
rect 2262 2459 2619 2501
rect -2175 2360 1979 2384
rect -2175 -2360 -2151 2360
rect 1955 -2360 1979 2360
rect -2175 -2384 1979 -2360
rect -258 -2716 62 -2384
rect 2262 -2459 2341 2459
rect 2577 -2459 2619 2459
rect 2262 -2501 2619 -2459
rect 2262 -2599 2582 -2501
rect 2262 -2641 2619 -2599
rect -2175 -2740 1979 -2716
rect -2175 -7460 -2151 -2740
rect 1955 -7460 1979 -2740
rect -2175 -7484 1979 -7460
rect -258 -7650 62 -7484
rect 2262 -7559 2341 -2641
rect 2577 -7559 2619 -2641
rect 2262 -7601 2619 -7559
rect 2262 -7650 2582 -7601
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2598 2600 2402 7600
string parameters w 24.0 l 24.0 val 1.17k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 87
string library sky130
<< end >>
