** sch_path: /home/hugodg/projects/temp-sensor/buffer/xschem/buffer_tb-dc.sch
**.subckt buffer_tb-dc
VIN1 in1 GND 1.2
.save i(vin1)
ibias vd ib 5u
VDD vd GND 1.8
.save i(vdd)
VSS vs GND 0
.save i(vss)
Cl out GND 4p m=1
X1 vd in1 out ib vs buffer-pex
**** begin user architecture code



.control
set color0=white
set color1=black

destroy all
save all
*dc ibias 0 20u 0.01u
dc VIN1 0.01 1.8 0.01
run
let err = abs(out-in1)
plot err ylabel 'Error (V)'
plot v(out) v(in1)


.endc

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /home/hugodg/projects/temp-sensor/buffer/xschem/buffer-pex.sym # of pins=5
** sym_path: /home/hugodg/projects/temp-sensor/buffer/xschem/buffer-pex.sym
** sch_path: /home/hugodg/projects/temp-sensor/buffer/xschem/buffer-pex.sch
.subckt buffer-pex vd in out ib gnd
*.iopin vd
*.iopin ib
*.iopin out
*.iopin in
*.iopin gnd
XM3 net2 net2 vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 out net4 gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 in net4 gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 net3 vd vd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 ib gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out net3 vd vd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out net1 gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net1 net2 vd vd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 net1 gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 ib ib gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


C0 net3 w_19600_3400# 0.0399f
C1 net3 in 1.06f
C2 net2 vd 2.85f
C3 a_14316_3522# vd 0.0215f
C4 a_19796_4422# vd 0.0104f
C5 gnd w_19600_3400# 0.0414f
C6 gnd in 0.0898f
C7 a_14316_4422# vd 0.0237f
C8 w_19600_3400# vd 0.0714f
C9 vd in 0.16f
C10 w_14120_3400# vd 0.116f
C11 w_19600_4300# vd 0.0724f
C12 w_14120_4300# vd 0.123f
C13 net1 out 2.63f
C14 net4 out 2.41f
C15 net3 out 2.19f
C16 net4 net1 0.0315f
C17 net3 net1 0.16f
C18 net4 ib 0.0512f
C19 net3 net4 1.5f
C20 a_21636_2682# in 0.0102f
C21 gnd out 1.84f
C22 vd out 1.05f
C23 net1 gnd 4.77f
C24 net4 gnd 0.596f
C25 ib gnd 0.163f
C26 net1 vd 1.48f
C27 net3 gnd 0.387f
C28 a_15696_2770# a_15438_2770# 0.0212f
C29 net3 vd 2.15f
C30 a_19996_3619# a_19738_3619# 0.0212f
C31 a_14258_3619# a_14516_3619# 0.0212f
C32 gnd vd 0.264f
C33 a_15696_2770# in 0.0215f
C34 a_19996_4519# a_19738_4519# 0.0212f
C35 net2 in 0.615f
C36 a_15496_2682# in 0.102f
C37 a_19996_3619# w_19600_3400# 0.0649f
C38 a_21636_1802# out 0.0539f
C39 a_19738_3619# w_19600_3400# 0.0649f
C40 w_19600_3400# a_19796_3522# 0.395f
C41 w_14120_3400# a_14258_3619# 0.0649f
C42 w_14120_3400# a_14516_3619# 0.0649f
C43 a_14316_3522# in 0.01f
C44 a_14516_4519# a_14258_4519# 0.0212f
C45 a_14316_3522# w_14120_3400# 0.395f
C46 a_19996_4519# w_19600_4300# 0.0649f
C47 w_19600_4300# a_19738_4519# 0.0649f
C48 w_19600_4300# a_19796_4422# 0.395f
C49 a_14516_4519# w_14120_4300# 0.0649f
C50 a_14556_1802# ib 0.0355f
C51 w_14120_4300# a_14258_4519# 0.0649f
C52 w_19600_3400# in 0.0115f
C53 w_14120_3400# in 0.0401f
C54 a_14316_4422# w_14120_4300# 0.395f
C55 w_19600_4300# w_19600_3400# 0.0394f
C56 w_14120_3400# w_14120_4300# 0.0394f
C57 net2 out 2.04f
C58 a_14498_1890# a_14756_1890# 0.0212f
C59 a_19796_3522# out 0.0116f
C60 net2 net1 1.99f
C61 net4 net2 1.32f
C62 a_21578_2770# a_21836_2770# 0.0212f
C63 net3 net2 0.338f
C64 a_21578_1890# a_21836_1890# 0.0212f
C65 w_19600_3400# out 0.0264f
C66 in out 1.56f
C67 net3 a_19796_3522# 0.0141f
C68 net1 in 0.296f
C69 net4 in 2.43f
C70 net2 gnd 0.342f
C71 ib in 0.0824f
C72 a_21836_1890# 0 0.0875f
C73 a_21578_1890# 0 0.0875f
C74 a_21636_1802# 0 0.6f
C75 a_14756_1890# 0 0.0875f
C76 a_14498_1890# 0 0.0875f
C77 a_14556_1802# 0 0.607f
C78 a_21836_2770# 0 0.0875f
C79 a_21578_2770# 0 0.0875f
C80 a_21636_2682# 0 0.6f
C81 a_15696_2770# 0 0.0875f
C82 a_15438_2770# 0 0.0875f
C83 a_15496_2682# 0 0.607f
C84 a_19996_3619# 0 0.0223f
C85 a_19738_3619# 0 0.0223f
C86 a_19796_3522# 0 0.225f
C87 a_14516_3619# 0 0.0223f
C88 a_14258_3619# 0 0.0223f
C89 a_14316_3522# 0 0.226f
C90 a_19996_4519# 0 0.0223f
C91 a_19738_4519# 0 0.0223f
C92 a_19796_4422# 0 0.226f
C93 a_14516_4519# 0 0.0223f
C94 a_14258_4519# 0 0.0223f
C95 a_14316_4422# 0 0.226f
C96 w_19600_3400# 0 1.6f
C97 w_14120_3400# 0 1.6f
C98 w_19600_4300# 0 1.6f
C99 w_14120_4300# 0 1.6f
C100 net4 0 1.22f
C101 ib 0 2.02f
C102 vd 0 19.5f
C103 gnd 0 -0.969f
C104 net1 0 21.9f
C105 net2 0 4.04f
C106 net3 0 3.79f
C107 in 0 6.74f
C108 out 0 11.9f


**** end user architecture code
XCc out net1 sky130_fd_pr__cap_mim_m3_2 W=21 L=21 MF=1 m=1
.ends

.GLOBAL GND
.end
