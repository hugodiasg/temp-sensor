magic
tech sky130A
magscale 1 2
timestamp 1645799662
<< metal4 >>
rect -2379 6959 2379 7000
rect -2379 2441 2123 6959
rect 2359 2441 2379 6959
rect -2379 2400 2379 2441
rect -2379 2259 2379 2300
rect -2379 -2259 2123 2259
rect 2359 -2259 2379 2259
rect -2379 -2300 2379 -2259
rect -2379 -2441 2379 -2400
rect -2379 -6959 2123 -2441
rect 2359 -6959 2379 -2441
rect -2379 -7000 2379 -6959
<< via4 >>
rect 2123 2441 2359 6959
rect 2123 -2259 2359 2259
rect 2123 -6959 2359 -2441
<< mimcap2 >>
rect -2279 6860 2121 6900
rect -2279 2540 -1807 6860
rect 1649 2540 2121 6860
rect -2279 2500 2121 2540
rect -2279 2160 2121 2200
rect -2279 -2160 -1807 2160
rect 1649 -2160 2121 2160
rect -2279 -2200 2121 -2160
rect -2279 -2540 2121 -2500
rect -2279 -6860 -1807 -2540
rect 1649 -6860 2121 -2540
rect -2279 -6900 2121 -6860
<< mimcap2contact >>
rect -1807 2540 1649 6860
rect -1807 -2160 1649 2160
rect -1807 -6860 1649 -2540
<< metal5 >>
rect -239 6884 81 7050
rect 2081 6959 2401 7050
rect -1831 6860 1673 6884
rect -1831 2540 -1807 6860
rect 1649 2540 1673 6860
rect -1831 2516 1673 2540
rect -239 2184 81 2516
rect 2081 2441 2123 6959
rect 2359 2441 2401 6959
rect 2081 2259 2401 2441
rect -1831 2160 1673 2184
rect -1831 -2160 -1807 2160
rect 1649 -2160 1673 2160
rect -1831 -2184 1673 -2160
rect -239 -2516 81 -2184
rect 2081 -2259 2123 2259
rect 2359 -2259 2401 2259
rect 2081 -2441 2401 -2259
rect -1831 -2540 1673 -2516
rect -1831 -6860 -1807 -2540
rect 1649 -6860 1673 -2540
rect -1831 -6884 1673 -6860
rect -239 -7050 81 -6884
rect 2081 -6959 2123 -2441
rect 2359 -6959 2401 -2441
rect 2081 -7050 2401 -6959
<< properties >>
string FIXED_BBOX -2379 2400 2221 7000
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
