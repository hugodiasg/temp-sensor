magic
tech sky130A
magscale 1 2
timestamp 1646014094
<< metal4 >>
rect -2681 7865 2681 7906
rect -2681 2743 2425 7865
rect 2661 2743 2681 7865
rect -2681 2702 2681 2743
rect -2681 2561 2681 2602
rect -2681 -2561 2425 2561
rect 2661 -2561 2681 2561
rect -2681 -2602 2681 -2561
rect -2681 -2743 2681 -2702
rect -2681 -7865 2425 -2743
rect 2661 -7865 2681 -2743
rect -2681 -7906 2681 -7865
<< via4 >>
rect 2425 2743 2661 7865
rect 2425 -2561 2661 2561
rect 2425 -7865 2661 -2743
<< mimcap2 >>
rect -2581 7766 2423 7806
rect -2581 2842 -2049 7766
rect 1891 2842 2423 7766
rect -2581 2802 2423 2842
rect -2581 2462 2423 2502
rect -2581 -2462 -2049 2462
rect 1891 -2462 2423 2462
rect -2581 -2502 2423 -2462
rect -2581 -2842 2423 -2802
rect -2581 -7766 -2049 -2842
rect 1891 -7766 2423 -2842
rect -2581 -7806 2423 -7766
<< mimcap2contact >>
rect -2049 2842 1891 7766
rect -2049 -2462 1891 2462
rect -2049 -7766 1891 -2842
<< metal5 >>
rect -239 7790 81 7956
rect 2383 7865 2703 7956
rect -2073 7766 1915 7790
rect -2073 2842 -2049 7766
rect 1891 2842 1915 7766
rect -2073 2818 1915 2842
rect -239 2486 81 2818
rect 2383 2743 2425 7865
rect 2661 2743 2703 7865
rect 2383 2561 2703 2743
rect -2073 2462 1915 2486
rect -2073 -2462 -2049 2462
rect 1891 -2462 1915 2462
rect -2073 -2486 1915 -2462
rect -239 -2818 81 -2486
rect 2383 -2561 2425 2561
rect 2661 -2561 2703 2561
rect 2383 -2743 2703 -2561
rect -2073 -2842 1915 -2818
rect -2073 -7766 -2049 -2842
rect 1891 -7766 1915 -2842
rect -2073 -7790 1915 -7766
rect -239 -7956 81 -7790
rect 2383 -7865 2425 -2743
rect 2661 -7865 2703 -2743
rect 2383 -7956 2703 -7865
<< properties >>
string FIXED_BBOX -2681 2702 2523 7906
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.019 l 25.019 val 1.27k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
