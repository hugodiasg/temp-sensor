magic
tech sky130A
timestamp 1644598236
<< metal4 >>
rect 2800 4470 3200 8400
rect 2800 4120 2830 4470
rect 3180 4120 3200 4470
rect 2800 4100 3200 4120
<< via4 >>
rect 2830 4120 3180 4470
<< metal5 >>
rect 0 7600 8000 8000
rect 0 6900 7300 7300
rect 0 400 400 6900
rect 700 6200 6600 6600
rect 700 1100 1100 6200
rect 1400 5500 5900 5900
rect 1400 1800 1800 5500
rect 2100 4800 5200 5200
rect 2100 2500 2500 4800
rect 2800 4470 3200 4500
rect 2800 4120 2830 4470
rect 3180 4120 3200 4470
rect 2800 3200 3200 4120
rect 4800 3200 5200 4800
rect 2800 2800 5200 3200
rect 5500 2500 5900 5500
rect 2100 2100 5900 2500
rect 6200 1800 6600 6200
rect 1400 1400 6600 1800
rect 6900 1100 7300 6900
rect 700 700 7300 1100
rect 7600 400 8000 7600
rect 0 0 8000 400
<< end >>
