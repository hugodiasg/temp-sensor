magic
tech sky130A
magscale 1 2
timestamp 1644768462
<< metal4 >>
rect -2539 7439 2539 7480
rect -2539 2601 2283 7439
rect 2519 2601 2539 7439
rect -2539 2560 2539 2601
rect -2539 2419 2539 2460
rect -2539 -2419 2283 2419
rect 2519 -2419 2539 2419
rect -2539 -2460 2539 -2419
rect -2539 -2601 2539 -2560
rect -2539 -7439 2283 -2601
rect 2519 -7439 2539 -2601
rect -2539 -7480 2539 -7439
<< via4 >>
rect 2283 2601 2519 7439
rect 2283 -2419 2519 2419
rect 2283 -7439 2519 -2601
<< mimcap2 >>
rect -2439 7340 2281 7380
rect -2439 2700 -1935 7340
rect 1777 2700 2281 7340
rect -2439 2660 2281 2700
rect -2439 2320 2281 2360
rect -2439 -2320 -1935 2320
rect 1777 -2320 2281 2320
rect -2439 -2360 2281 -2320
rect -2439 -2700 2281 -2660
rect -2439 -7340 -1935 -2700
rect 1777 -7340 2281 -2700
rect -2439 -7380 2281 -7340
<< mimcap2contact >>
rect -1935 2700 1777 7340
rect -1935 -2320 1777 2320
rect -1935 -7340 1777 -2700
<< metal5 >>
rect -239 7364 81 7530
rect 2241 7439 2561 7530
rect -1959 7340 1801 7364
rect -1959 2700 -1935 7340
rect 1777 2700 1801 7340
rect -1959 2676 1801 2700
rect -239 2344 81 2676
rect 2241 2601 2283 7439
rect 2519 2601 2561 7439
rect 2241 2419 2561 2601
rect -1959 2320 1801 2344
rect -1959 -2320 -1935 2320
rect 1777 -2320 1801 2320
rect -1959 -2344 1801 -2320
rect -239 -2676 81 -2344
rect 2241 -2419 2283 2419
rect 2519 -2419 2561 2419
rect 2241 -2601 2561 -2419
rect -1959 -2700 1801 -2676
rect -1959 -7340 -1935 -2700
rect 1777 -7340 1801 -2700
rect -1959 -7364 1801 -7340
rect -239 -7530 81 -7364
rect 2241 -7439 2283 -2601
rect 2519 -7439 2561 -2601
rect 2241 -7530 2561 -7439
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2539 2560 2381 7480
string parameters w 23.6 l 23.6 val 1.131k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
