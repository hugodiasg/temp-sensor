magic
tech sky130A
magscale 1 2
timestamp 1644355690
<< pwell >>
rect -1436 -654 1436 654
<< psubdiff >>
rect -1400 584 -1304 618
rect 1304 584 1400 618
rect -1400 522 -1366 584
rect 1366 522 1400 584
rect -1400 -584 -1366 -522
rect 1366 -584 1400 -522
rect -1400 -618 -1304 -584
rect 1304 -618 1400 -584
<< psubdiffcont >>
rect -1304 584 1304 618
rect -1400 -522 -1366 522
rect 1366 -522 1400 522
rect -1304 -618 1304 -584
<< xpolycontact >>
rect -1270 56 -124 488
rect -1270 -488 -124 -56
rect 124 56 1270 488
rect 124 -488 1270 -56
<< ppolyres >>
rect -1270 -56 -124 56
rect 124 -56 1270 56
<< locali >>
rect -1400 584 -1304 618
rect 1304 584 1400 618
rect -1400 522 -1366 584
rect -1400 -584 -1366 -522
rect -1400 -618 -1304 -584
rect 1304 -618 1400 -584
<< viali >>
rect 1366 522 1400 584
rect -1254 73 -140 470
rect 140 73 1254 470
rect -1254 -470 -140 -73
rect 140 -470 1254 -73
rect 1366 -522 1400 522
rect 1366 -584 1400 -522
<< metal1 >>
rect 1360 584 1406 596
rect -1266 470 -128 476
rect -1266 73 -1254 470
rect -140 73 -128 470
rect -1266 67 -128 73
rect 128 470 1266 476
rect 128 73 140 470
rect 1254 73 1266 470
rect 128 67 1266 73
rect -1266 -73 -128 -67
rect -1266 -470 -1254 -73
rect -140 -470 -128 -73
rect -1266 -476 -128 -470
rect 128 -73 1266 -67
rect 128 -470 140 -73
rect 1254 -470 1266 -73
rect 128 -476 1266 -470
rect 1360 -584 1366 584
rect 1400 -584 1406 584
rect 1360 -596 1406 -584
<< res5p73 >>
rect -1272 -58 -122 58
rect 122 -58 1272 58
<< properties >>
string gencell sky130_fd_pr__res_high_po_5p73
string FIXED_BBOX -1383 -601 1383 601
string parameters w 5.730 l 0.56 m 1 nx 2 wmin 5.730 lmin 0.50 rho 319.8 val 37.951 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 100
string library sky130
<< end >>
