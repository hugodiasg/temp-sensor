* NGSPICE file created from ask-modulator.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_NVRUDW w_n201_n1098# a_n35_500# a_n35_n932#
X0 a_n35_n932# a_n35_500# w_n201_n1098# sky130_fd_pr__res_xhigh_po_0p35 l=5e+06u
C0 a_n35_n932# w_n201_n1098# 1.08fF
C1 a_n35_500# w_n201_n1098# 1.08fF
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ML7W5H a_n108_n870# a_n50_n958# w_n278_n1128#
+ a_50_n870#
X0 a_50_n870# a_n50_n958# a_n108_n870# w_n278_n1128# sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=8.7e+06u l=500000u
C0 a_50_n870# a_n108_n870# 1.16fF
C1 a_50_n870# w_n278_n1128# 0.87fF
C2 a_n108_n870# w_n278_n1128# 0.87fF
C3 a_n50_n958# w_n278_n1128# 0.52fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_QKF9RA c2_n2379_n7200# m4_n2479_n7300# VSUBS
X0 c2_n2379_n7200# m4_n2479_n7300# sky130_fd_pr__cap_mim_m3_2 l=2.3e+07u w=2.3e+07u
X1 c2_n2379_n7200# m4_n2479_n7300# sky130_fd_pr__cap_mim_m3_2 l=2.3e+07u w=2.3e+07u
X2 c2_n2379_n7200# m4_n2479_n7300# sky130_fd_pr__cap_mim_m3_2 l=2.3e+07u w=2.3e+07u
C0 m4_n2479_n7300# c2_n2379_n7200# 106.47fF
C1 c2_n2379_n7200# VSUBS 0.26fF
C2 m4_n2479_n7300# VSUBS 28.22fF
.ends

.subckt ask-modulator in out gnd
XXR1 gnd out out sky130_fd_pr__res_xhigh_po_0p35_NVRUDW
XXM1 gnd in gnd out sky130_fd_pr__nfet_g5v0d10v5_ML7W5H
XXC0 out out gnd sky130_fd_pr__cap_mim_m3_2_QKF9RA
X0 out out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
X1 out in.t0 gnd gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=0u l=0u
X2 out out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
X3 out out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 gnd.n0 gnd 0.619
R1 gnd gnd.n0 0.07
R2 gnd.n0 gnd 0.062
R3 in in.t0 446.385
C0 out in 0.05fF
C1 out gnd 323.51fF
C2 in gnd 1.10fF
.ends

