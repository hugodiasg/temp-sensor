magic
tech sky130A
magscale 1 2
timestamp 1645139004
<< mvpsubdiff >>
rect -23398 -19130 -23374 -17659
rect -21874 -19130 -21850 -17659
<< mvpsubdiffcont >>
rect -23374 -19130 -21874 -17659
<< locali >>
rect -23390 -19130 -23374 -17659
rect -21874 -19130 -21858 -17659
<< viali >>
rect -23186 -17806 -22020 -17799
rect -23205 -19005 -21999 -17806
<< metal1 >>
rect -24800 11200 -21400 11400
rect -24800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -24800 9800 -21400 10000
rect 9600 -7200 11400 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11400 -7200
rect 9600 -8400 11400 -8200
rect -24800 -17799 -21800 -17600
rect -24800 -17800 -23186 -17799
rect -22020 -17800 -21800 -17799
rect -24800 -17806 -23200 -17800
rect -22000 -17806 -21800 -17800
rect -24800 -19005 -23205 -17806
rect -21999 -19005 -21800 -17806
rect -24800 -19200 -21800 -19005
<< via1 >>
rect -22600 10000 -21600 11200
rect 9800 -8200 10800 -7200
rect -23200 -17806 -23186 -17800
rect -23186 -17806 -22020 -17800
rect -22020 -17806 -22000 -17800
rect -23200 -19000 -22000 -17806
<< metal2 >>
rect -22800 11200 -21400 11400
rect -22800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -22800 9800 -21400 10000
rect 9600 -7200 11000 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect 9600 -8400 11000 -8200
rect -23400 -17800 -21800 -17600
rect -23400 -19000 -23200 -17800
rect -22000 -19000 -21800 -17800
rect -23400 -19200 -21800 -19000
<< via2 >>
rect -22600 10000 -21600 11200
rect 9800 -8200 10800 -7200
rect -23200 -19000 -22000 -17800
<< metal3 >>
rect -22800 11200 -21400 11400
rect -22800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -22800 9800 -21400 10000
rect 9600 -7200 11000 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect 9600 -8400 11000 -8200
rect -23400 -17800 -21800 -17600
rect -23400 -19000 -23200 -17800
rect -22000 -19000 -21800 -17800
rect -23400 -19200 -21800 -19000
<< via3 >>
rect -22600 10000 -21600 11200
rect 9800 -8200 10800 -7200
rect -23200 -19000 -22000 -17800
<< metal4 >>
rect -22800 11200 -21400 11400
rect -22800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -22800 9800 -21400 10000
rect -24600 7049 -19962 7090
rect -24600 2651 -20218 7049
rect -19982 2651 -19962 7049
rect -24600 2610 -19962 2651
rect -19400 7049 -14762 7090
rect -19400 2651 -15018 7049
rect -14782 2651 -14762 7049
rect -19400 2610 -14762 2651
rect -14000 7049 -9362 7090
rect -14000 2651 -9618 7049
rect -9382 2651 -9362 7049
rect -14000 2610 -9362 2651
rect -24600 2469 -19962 2510
rect -24600 -1929 -20218 2469
rect -19982 -1929 -19962 2469
rect -24600 -1970 -19962 -1929
rect -19400 2469 -14762 2510
rect -19400 -1929 -15018 2469
rect -14782 -1929 -14762 2469
rect -19400 -1970 -14762 -1929
rect -14000 2469 -9362 2510
rect -14000 -1929 -9618 2469
rect -9382 -1929 -9362 2469
rect -14000 -1970 -9362 -1929
rect -24600 -2111 -19962 -2070
rect -24600 -6509 -20218 -2111
rect -19982 -6509 -19962 -2111
rect -24600 -6550 -19962 -6509
rect -19400 -2111 -14762 -2070
rect -19400 -6509 -15018 -2111
rect -14782 -6509 -14762 -2111
rect -19400 -6550 -14762 -6509
rect -14000 -2111 -9362 -2070
rect -14000 -6509 -9618 -2111
rect -9382 -6509 -9362 -2111
rect -14000 -6550 -9362 -6509
rect -23000 -8200 -21600 -6550
rect -17600 -8200 -16200 -6550
rect -11800 -8200 -10400 -6550
rect 2680 -7000 4360 1998
rect -23000 -9600 -10400 -8200
rect 2600 -7200 4400 -7000
rect 2600 -8200 2800 -7200
rect 4200 -8200 4400 -7200
rect 2600 -8400 4400 -8200
rect 9600 -7200 11000 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect 9600 -8400 11000 -8200
rect -23000 -17600 -21600 -9600
rect -11000 -10407 -5314 -10366
rect -11000 -15853 -5570 -10407
rect -5334 -15853 -5314 -10407
rect -11000 -15894 -5314 -15853
rect -4800 -10407 886 -10366
rect -4800 -15853 630 -10407
rect 866 -15853 886 -10407
rect -4800 -15894 886 -15853
rect 1200 -10407 6886 -10366
rect 1200 -15853 6630 -10407
rect 6866 -15853 6886 -10407
rect 1200 -15894 6886 -15853
rect 7600 -10407 13286 -10366
rect 7600 -15853 13030 -10407
rect 13266 -15853 13286 -10407
rect 7600 -15894 13286 -15853
rect -23425 -17800 -21600 -17600
rect -23425 -19000 -23200 -17800
rect -22000 -19000 -21600 -17800
rect -23425 -19233 -21600 -19000
rect -23000 -28200 -21600 -19233
rect -11000 -16035 -5314 -15994
rect -11000 -21481 -5570 -16035
rect -5334 -21481 -5314 -16035
rect -11000 -21522 -5314 -21481
rect -4800 -16035 886 -15994
rect -4800 -21481 630 -16035
rect 866 -21481 886 -16035
rect -4800 -21522 886 -21481
rect 1200 -16035 6886 -15994
rect 1200 -21481 6630 -16035
rect 6866 -21481 6886 -16035
rect 1200 -21522 6886 -21481
rect 7600 -16035 13286 -15994
rect 7600 -21481 13030 -16035
rect 13266 -21481 13286 -16035
rect 7600 -21522 13286 -21481
rect -11000 -21663 -5314 -21622
rect -11000 -27109 -5570 -21663
rect -5334 -27109 -5314 -21663
rect -11000 -27150 -5314 -27109
rect -4800 -21663 886 -21622
rect -4800 -27109 630 -21663
rect 866 -27109 886 -21663
rect -4800 -27150 886 -27109
rect 1200 -21663 6886 -21622
rect 1200 -27109 6630 -21663
rect 6866 -27109 6886 -21663
rect 1200 -27150 6886 -27109
rect 7600 -21663 13286 -21622
rect 7600 -27109 13030 -21663
rect 13266 -27109 13286 -21663
rect 7600 -27150 13286 -27109
rect -9000 -28200 -7400 -27150
rect -23000 -28400 -7400 -28200
rect -3400 -28400 -1800 -27150
rect 3400 -28400 5000 -27150
rect 9600 -28400 11200 -27150
rect -23000 -29800 11200 -28400
<< via4 >>
rect -22600 10000 -21600 11200
rect -20218 2651 -19982 7049
rect -15018 2651 -14782 7049
rect -9618 2651 -9382 7049
rect -20218 -1929 -19982 2469
rect -15018 -1929 -14782 2469
rect -9618 -1929 -9382 2469
rect -20218 -6509 -19982 -2111
rect -15018 -6509 -14782 -2111
rect -9618 -6509 -9382 -2111
rect 2800 -8200 4200 -7200
rect 9800 -8200 10800 -7200
rect -5570 -15853 -5334 -10407
rect 630 -15853 866 -10407
rect 6630 -15853 6866 -10407
rect 13030 -15853 13266 -10407
rect -5570 -21481 -5334 -16035
rect 630 -21481 866 -16035
rect 6630 -21481 6866 -16035
rect 13030 -21481 13266 -16035
rect -5570 -27109 -5334 -21663
rect 630 -27109 866 -21663
rect 6630 -27109 6866 -21663
rect 13030 -27109 13266 -21663
<< mimcap2 >>
rect -24500 6950 -20220 6990
rect -24500 2750 -24040 6950
rect -20680 2750 -20220 6950
rect -24500 2710 -20220 2750
rect -19300 6950 -15020 6990
rect -19300 2750 -18840 6950
rect -15480 2750 -15020 6950
rect -19300 2710 -15020 2750
rect -13900 6950 -9620 6990
rect -13900 2750 -13440 6950
rect -10080 2750 -9620 6950
rect -13900 2710 -9620 2750
rect -24500 2370 -20220 2410
rect -24500 -1830 -24040 2370
rect -20680 -1830 -20220 2370
rect -24500 -1870 -20220 -1830
rect -19300 2370 -15020 2410
rect -19300 -1830 -18840 2370
rect -15480 -1830 -15020 2370
rect -19300 -1870 -15020 -1830
rect -13900 2370 -9620 2410
rect -13900 -1830 -13440 2370
rect -10080 -1830 -9620 2370
rect -13900 -1870 -9620 -1830
rect -24500 -2210 -20220 -2170
rect -24500 -6410 -24040 -2210
rect -20680 -6410 -20220 -2210
rect -24500 -6450 -20220 -6410
rect -19300 -2210 -15020 -2170
rect -19300 -6410 -18840 -2210
rect -15480 -6410 -15020 -2210
rect -19300 -6450 -15020 -6410
rect -13900 -2210 -9620 -2170
rect -13900 -6410 -13440 -2210
rect -10080 -6410 -9620 -2210
rect -13900 -6450 -9620 -6410
rect -10900 -10506 -5572 -10466
rect -10900 -15754 -10335 -10506
rect -6137 -15754 -5572 -10506
rect -10900 -15794 -5572 -15754
rect -4700 -10506 628 -10466
rect -4700 -15754 -4135 -10506
rect 63 -15754 628 -10506
rect -4700 -15794 628 -15754
rect 1300 -10506 6628 -10466
rect 1300 -15754 1865 -10506
rect 6063 -15754 6628 -10506
rect 1300 -15794 6628 -15754
rect 7700 -10506 13028 -10466
rect 7700 -15754 8265 -10506
rect 12463 -15754 13028 -10506
rect 7700 -15794 13028 -15754
rect -10900 -16134 -5572 -16094
rect -10900 -21382 -10335 -16134
rect -6137 -21382 -5572 -16134
rect -10900 -21422 -5572 -21382
rect -4700 -16134 628 -16094
rect -4700 -21382 -4135 -16134
rect 63 -21382 628 -16134
rect -4700 -21422 628 -21382
rect 1300 -16134 6628 -16094
rect 1300 -21382 1865 -16134
rect 6063 -21382 6628 -16134
rect 1300 -21422 6628 -21382
rect 7700 -16134 13028 -16094
rect 7700 -21382 8265 -16134
rect 12463 -21382 13028 -16134
rect 7700 -21422 13028 -21382
rect -10900 -21762 -5572 -21722
rect -10900 -27010 -10335 -21762
rect -6137 -27010 -5572 -21762
rect -10900 -27050 -5572 -27010
rect -4700 -21762 628 -21722
rect -4700 -27010 -4135 -21762
rect 63 -27010 628 -21762
rect -4700 -27050 628 -27010
rect 1300 -21762 6628 -21722
rect 1300 -27010 1865 -21762
rect 6063 -27010 6628 -21762
rect 1300 -27050 6628 -27010
rect 7700 -21762 13028 -21722
rect 7700 -27010 8265 -21762
rect 12463 -27010 13028 -21762
rect 7700 -27050 13028 -27010
<< mimcap2contact >>
rect -24040 2750 -20680 6950
rect -18840 2750 -15480 6950
rect -13440 2750 -10080 6950
rect -24040 -1830 -20680 2370
rect -18840 -1830 -15480 2370
rect -13440 -1830 -10080 2370
rect -24040 -6410 -20680 -2210
rect -18840 -6410 -15480 -2210
rect -13440 -6410 -10080 -2210
rect -10335 -15754 -6137 -10506
rect -4135 -15754 63 -10506
rect 1865 -15754 6063 -10506
rect 8265 -15754 12463 -10506
rect -10335 -21382 -6137 -16134
rect -4135 -21382 63 -16134
rect 1865 -21382 6063 -16134
rect 8265 -21382 12463 -16134
rect -10335 -27010 -6137 -21762
rect -4135 -27010 63 -21762
rect 1865 -27010 6063 -21762
rect 8265 -27010 12463 -21762
<< metal5 >>
rect -22840 11200 11200 11480
rect -22840 10000 -22600 11200
rect -21600 10000 11200 11200
rect -22840 9800 11200 10000
rect -22800 6974 -21400 9800
rect -20260 7049 -19940 7140
rect -24064 6950 -20656 6974
rect -24064 2750 -24040 6950
rect -20680 2750 -20656 6950
rect -24064 2726 -20656 2750
rect -22520 2394 -22200 2726
rect -20260 2651 -20218 7049
rect -19982 2651 -19940 7049
rect -17600 6974 -16200 9800
rect -11800 7140 -10200 9800
rect -6800 7520 8920 9200
rect -15060 7049 -14740 7140
rect -18864 6950 -15456 6974
rect -18864 2750 -18840 6950
rect -15480 2750 -15456 6950
rect -18864 2726 -15456 2750
rect -20260 2469 -19940 2651
rect -24064 2370 -20656 2394
rect -24064 -1830 -24040 2370
rect -20680 -1830 -20656 2370
rect -24064 -1854 -20656 -1830
rect -22520 -2186 -22200 -1854
rect -20260 -1929 -20218 2469
rect -19982 -1929 -19940 2469
rect -17320 2394 -17000 2726
rect -15060 2651 -15018 7049
rect -14782 2651 -14740 7049
rect -11920 6974 -10200 7140
rect -9660 7049 -9340 7140
rect -13464 6950 -10056 6974
rect -13464 2750 -13440 6950
rect -10080 2750 -10056 6950
rect -13464 2726 -10056 2750
rect -15060 2469 -14740 2651
rect -18864 2370 -15456 2394
rect -18864 -1830 -18840 2370
rect -15480 -1830 -15456 2370
rect -18864 -1854 -15456 -1830
rect -20260 -2111 -19940 -1929
rect -24064 -2210 -20656 -2186
rect -24064 -6410 -24040 -2210
rect -20680 -6410 -20656 -2210
rect -24064 -6434 -20656 -6410
rect -22520 -6600 -22200 -6434
rect -20260 -6509 -20218 -2111
rect -19982 -6509 -19940 -2111
rect -17320 -2186 -17000 -1854
rect -15060 -1929 -15018 2469
rect -14782 -1929 -14740 2469
rect -11920 2394 -11600 2726
rect -9660 2651 -9618 7049
rect -9382 2651 -9340 7049
rect -9660 2469 -9340 2651
rect -13464 2370 -10056 2394
rect -13464 -1830 -13440 2370
rect -10080 -1830 -10056 2370
rect -13464 -1854 -10056 -1830
rect -15060 -2111 -14740 -1929
rect -18864 -2210 -15456 -2186
rect -18864 -6410 -18840 -2210
rect -15480 -6410 -15456 -2210
rect -18864 -6434 -15456 -6410
rect -20260 -6600 -19940 -6509
rect -17320 -6600 -17000 -6434
rect -15060 -6509 -15018 -2111
rect -14782 -6509 -14740 -2111
rect -11920 -2186 -11600 -1854
rect -9660 -1929 -9618 2469
rect -9382 -1929 -9340 2469
rect -9660 -2111 -9340 -1929
rect -13464 -2210 -10056 -2186
rect -13464 -6410 -13440 -2210
rect -10080 -6410 -10056 -2210
rect -13464 -6434 -10056 -6410
rect -15060 -6600 -14740 -6509
rect -11920 -6600 -11600 -6434
rect -9660 -6509 -9618 -2111
rect -9382 -6509 -9340 -2111
rect -9660 -6600 -9340 -6509
rect -6800 -4842 -5122 7520
rect -4522 5240 6640 6920
rect -4522 -2562 -2842 5240
rect -2242 2960 4360 4640
rect -2242 -282 -562 2960
rect 2680 318 4360 2960
rect 4960 -282 6640 5240
rect -2242 -1962 6640 -282
rect 7240 -2562 8920 7520
rect -4522 -4242 8920 -2562
rect 9520 -4842 11200 9800
rect -6800 -6520 11200 -4842
rect -8800 -7200 11000 -7000
rect -8800 -8200 2800 -7200
rect 4200 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect -8800 -8400 11000 -8200
rect -8800 -10482 -7600 -8400
rect -5612 -10407 -5292 -10316
rect -10359 -10506 -6113 -10482
rect -10359 -15754 -10335 -10506
rect -6137 -15754 -6113 -10506
rect -10359 -15778 -6113 -15754
rect -8396 -16110 -8076 -15778
rect -5612 -15853 -5570 -10407
rect -5334 -15853 -5292 -10407
rect -2600 -10482 -1400 -8400
rect 588 -10407 908 -10316
rect -4159 -10506 87 -10482
rect -4159 -15754 -4135 -10506
rect 63 -15754 87 -10506
rect -4159 -15778 87 -15754
rect -5612 -16035 -5292 -15853
rect -10359 -16134 -6113 -16110
rect -10359 -21382 -10335 -16134
rect -6137 -21382 -6113 -16134
rect -10359 -21406 -6113 -21382
rect -8396 -21738 -8076 -21406
rect -5612 -21481 -5570 -16035
rect -5334 -21481 -5292 -16035
rect -2196 -16110 -1876 -15778
rect 588 -15853 630 -10407
rect 866 -15853 908 -10407
rect 3600 -10482 4800 -8400
rect 6588 -10407 6908 -10316
rect 1841 -10506 6087 -10482
rect 1841 -15754 1865 -10506
rect 6063 -15754 6087 -10506
rect 1841 -15778 6087 -15754
rect 588 -16035 908 -15853
rect -4159 -16134 87 -16110
rect -4159 -21382 -4135 -16134
rect 63 -21382 87 -16134
rect -4159 -21406 87 -21382
rect -5612 -21663 -5292 -21481
rect -10359 -21762 -6113 -21738
rect -10359 -27010 -10335 -21762
rect -6137 -27010 -6113 -21762
rect -10359 -27034 -6113 -27010
rect -8396 -27200 -8076 -27034
rect -5612 -27109 -5570 -21663
rect -5334 -27109 -5292 -21663
rect -2196 -21738 -1876 -21406
rect 588 -21481 630 -16035
rect 866 -21481 908 -16035
rect 3804 -16110 4124 -15778
rect 6588 -15853 6630 -10407
rect 6866 -15853 6908 -10407
rect 9800 -10482 11000 -8400
rect 12988 -10407 13308 -10316
rect 8241 -10506 12487 -10482
rect 8241 -15754 8265 -10506
rect 12463 -15754 12487 -10506
rect 8241 -15778 12487 -15754
rect 6588 -16035 6908 -15853
rect 1841 -16134 6087 -16110
rect 1841 -21382 1865 -16134
rect 6063 -21382 6087 -16134
rect 1841 -21406 6087 -21382
rect 588 -21663 908 -21481
rect -4159 -21762 87 -21738
rect -4159 -27010 -4135 -21762
rect 63 -27010 87 -21762
rect -4159 -27034 87 -27010
rect -5612 -27200 -5292 -27109
rect -2196 -27200 -1876 -27034
rect 588 -27109 630 -21663
rect 866 -27109 908 -21663
rect 3804 -21738 4124 -21406
rect 6588 -21481 6630 -16035
rect 6866 -21481 6908 -16035
rect 10204 -16110 10524 -15778
rect 12988 -15853 13030 -10407
rect 13266 -15853 13308 -10407
rect 12988 -16035 13308 -15853
rect 8241 -16134 12487 -16110
rect 8241 -21382 8265 -16134
rect 12463 -21382 12487 -16134
rect 8241 -21406 12487 -21382
rect 6588 -21663 6908 -21481
rect 1841 -21762 6087 -21738
rect 1841 -27010 1865 -21762
rect 6063 -27010 6087 -21762
rect 1841 -27034 6087 -27010
rect 588 -27200 908 -27109
rect 3804 -27200 4124 -27034
rect 6588 -27109 6630 -21663
rect 6866 -27109 6908 -21663
rect 10204 -21738 10524 -21406
rect 12988 -21481 13030 -16035
rect 13266 -21481 13308 -16035
rect 12988 -21663 13308 -21481
rect 8241 -21762 12487 -21738
rect 8241 -27010 8265 -21762
rect 12463 -27010 12487 -21762
rect 8241 -27034 12487 -27010
rect 6588 -27200 6908 -27109
rect 10204 -27200 10524 -27034
rect 12988 -27109 13030 -21663
rect 13266 -27109 13308 -21663
rect 12988 -27200 13308 -27109
<< labels >>
flabel metal1 11200 -8000 11400 -7800 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 -24800 10400 -24600 10600 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 -24800 -18400 -24600 -18200 0 FreeSans 256 0 0 0 gnd
port 0 nsew
<< end >>
