* NGSPICE file created from device-complete.ext - technology: sky130A

.subckt device-complete gnd clk out_sigma vts ib out_buff vd out vpwr
X0 gnd.t71 buffer_0.d out_buff.t5 gnd.t70 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 a_16688_5320# a_16854_3988# gnd.t91 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X2 vd.t68 buffer_0.a.t17 buffer_0.d vd.t67 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 sensor_0.a.t11 sensor_0.b.t20 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 out_buff.t2 buffer_0.d gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 sensor_0.b.t16 sensor_0.b.t15 gnd.t72 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 a_15868_2881# a_14791_2515# a_15706_2515# vpwr.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 gnd.t130 vpwr.t30 a_15403_2515# gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_15546_5320# a_15712_3988# gnd.t16 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X9 vd.t66 buffer_0.a.t18 buffer_0.d vd.t65 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X10 buffer_0.a.t16 buffer_0.a.t14 buffer_0.a.t15 gnd.t164 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X11 gnd.t154 sensor_0.b.t21 vtd.t7 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X12 a_15141_2515# a_14791_2515# a_15046_2515# vpwr.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X13 sensor_0.c sensor_0.c sensor_0.c vd.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=1
X14 buffer_0.c.t20 vts.t25 buffer_0.b.t3 gnd.t140 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X15 gnd.t118 gnd.t116 gnd.t117 gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X16 a_14550_5320# a_14716_3988# gnd.t9 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X17 a_15815_2515# a_14625_2515# a_15706_2515# gnd.t29 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X18 vd.t64 buffer_0.a.t19 buffer_0.d vd.t63 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X19 buffer_0.c.t9 out_buff.t21 buffer_0.a.t9 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 gnd.t165 sensor_0.b.t13 sensor_0.b.t14 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X21 vts.t16 vtd.t20 vtd.t21 vts.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X22 a_16356_5320# a_16522_3988# gnd.t8 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X23 vd.t23 vd.t21 vd.t23 vd.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X24 buffer_0.c.t19 vts.t26 buffer_0.b.t0 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X25 gnd.t160 ib.t0 ib.t1 gnd.t159 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 buffer_0.d buffer_0.d gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 gnd.t115 gnd.t113 gnd.t114 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X28 vtd.t13 vtd.t12 vts.t14 vts.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 gnd.t14 sensor_0.b.t22 sensor_0.a.t10 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X30 vd.t30 buffer_0.b.t10 out_buff.t14 vd.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X31 gnd.t112 gnd.t110 gnd.t111 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X32 vtd.t6 sensor_0.b.t23 gnd.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X33 out_sigma.t0 a_16445_2515# vpwr.t29 vpwr.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X34 gnd.t65 buffer_0.d out_buff.t8 gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 vts.t12 vtd.t14 vtd.t15 vts.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 buffer_0.c.t8 out_buff.t22 buffer_0.a.t8 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 vtd.t5 sensor_0.b.t24 gnd.t92 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X38 vpwr.t7 clk.t0 a_14625_2515# vpwr.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X39 out_buff.t11 buffer_0.d gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X40 a_17020_5320# sigma-delta_0.x1.Q gnd.t23 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X41 a_15237_2515# a_14791_2515# a_15141_2515# gnd.t134 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X42 a_15706_2515# a_14625_2515# a_15359_2757# vpwr.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X43 vtd.t17 vtd.t16 vts.t10 vts.t9 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X44 vd.t80 a_6126_29386# gnd.t168 sky130_fd_pr__res_xhigh_po_0p35 l=5
X45 sensor_0.b.t19 vtd.t24 sensor_0.c vd.t39 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X46 a_15359_2757# a_15141_2515# vpwr.t11 vpwr.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X47 gnd.t25 clk.t1 a_14625_2515# gnd.t24 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X48 buffer_0.a.t11 buffer_0.a.t10 vd.t62 vd.t61 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X49 gnd.t75 sensor_0.b.t11 sensor_0.b.t12 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X50 vpwr.t9 a_15706_2515# a_15881_2489# vpwr.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X51 vts.t8 vtd.t18 vtd.t19 vts.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X52 a_15046_2515# sigma-delta_0.x1.D vpwr.t27 vpwr.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X53 vd.t41 sensor_0.a.t2 sensor_0.a.t3 vd.t40 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X54 gnd.t61 buffer_0.d buffer_0.d gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X55 a_15881_2489# a_15706_2515# a_16060_2515# gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X56 buffer_0.a.t2 out_buff.t23 buffer_0.c.t7 gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X57 sensor_0.b.t10 sensor_0.b.t9 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X58 a_14882_5320# a_15048_3988# gnd.t12 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X59 buffer_0.d buffer_0.a.t20 vd.t60 vd.t59 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X60 gnd.t85 sensor_0.b.t25 sensor_0.a.t9 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X61 buffer_0.c.t18 vts.t27 buffer_0.b.t5 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X62 buffer_0.c.t17 vts.t28 buffer_0.b.t4 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X63 buffer_0.b.t1 vts.t29 buffer_0.c.t16 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X64 buffer_0.b.t7 vts.t30 buffer_0.c.t15 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X65 sigma-delta_0.x1.Q a_15881_2489# gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X66 vd.t58 buffer_0.a.t21 buffer_0.d vd.t57 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X67 buffer_0.c.t10 ib.t5 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X68 vts.t24 vts.t21 vts.t23 vts.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X69 buffer_0.c.t6 out_buff.t24 buffer_0.a.t1 gnd.t125 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X70 gnd.t59 buffer_0.d buffer_0.d gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X71 gnd.t57 buffer_0.d buffer_0.d gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X72 a_15359_2757# a_15141_2515# gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X73 vpwr.t17 a_15359_2757# a_15249_2881# vpwr.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X74 buffer_0.d buffer_0.a.t22 vd.t56 vd.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X75 a_15706_2515# a_14791_2515# a_15359_2757# gnd.t133 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X76 gnd.t90 sensor_0.b.t26 vtd.t4 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X77 vd.t70 vtd.t25 vts.t6 vd.t69 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X78 vd.t54 buffer_0.a.t23 buffer_0.d vd.t53 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X79 a_15214_5320# a_15380_3988# gnd.t11 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X80 vd.t20 vd.t17 vd.t19 vd.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X81 buffer_0.d buffer_0.a.t24 vd.t52 vd.t51 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X82 buffer_0.a.t13 buffer_0.a.t12 buffer_0.a.t13 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X83 gnd.t109 gnd.t107 gnd.t108 gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X84 sensor_0.c vtd.t26 sensor_0.b.t18 vd.t36 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X85 buffer_0.a.t5 out_buff.t25 buffer_0.c.t5 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X86 out_sigma.t1 a_16445_2515# gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X87 buffer_0.d buffer_0.d gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X88 sensor_0.a.t8 sensor_0.b.t27 gnd.t89 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X89 sensor_0.a.t7 sensor_0.b.t28 gnd.t166 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X90 sigma-delta_0.x1.Q a_15881_2489# vpwr.t23 vpwr.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.213 ps=1.67 w=1 l=0.15
X91 sensor_0.a.t1 sensor_0.a.t0 vd.t74 vd.t73 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X92 gnd.t53 buffer_0.d out_buff.t4 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X93 vd.t83 out.t3 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X94 a_16060_2515# vpwr.t31 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X95 vd.t16 vd.t13 vd.t15 vd.t14 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X96 out_buff.t10 buffer_0.d gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X97 a_16024_5320# a_16190_3988# gnd.t135 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X98 sensor_0.b.t8 sensor_0.b.t7 gnd.t147 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X99 gnd.t4 sensor_0.b.t29 vtd.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X100 vd.t28 buffer_0.b.t11 out_buff.t13 vd.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X101 a_16688_5320# a_16522_3988# gnd.t162 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X102 vd.t12 vd.t9 vd.t11 vd.t10 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X103 buffer_0.a.t6 out_buff.t26 buffer_0.c.t4 gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X104 sensor_0.c sensor_0.a.t12 sensor_0.d vd.t75 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X105 sensor_0.d sensor_0.a.t13 sensor_0.c vd.t78 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X106 a_15546_5320# a_15380_3988# gnd.t153 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X107 vpwr.t21 a_15881_2489# a_15868_2881# vpwr.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X108 buffer_0.c.t3 out_buff.t27 buffer_0.a.t0 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X109 gnd.t106 gnd.t104 gnd.t105 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X110 gnd.t103 gnd.t101 gnd.t102 gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X111 gnd.t100 gnd.t97 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X112 vd.t8 vd.t5 vd.t7 vd.t6 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X113 buffer_0.d buffer_0.d gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X114 a_15046_2515# sigma-delta_0.x1.D gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X115 gnd.t138 sensor_0.b.t5 sensor_0.b.t6 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X116 vtd.t11 vtd.t10 vts.t5 vts.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X117 vd.t38 buffer_0.b.t12 out_buff.t16 vd.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X118 gnd.t47 buffer_0.d out_buff.t7 gnd.t46 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X119 gnd.t45 buffer_0.d out_buff.t6 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X120 gnd.t88 sensor_0.b.t30 sensor_0.a.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X121 a_15141_2515# a_14625_2515# a_15046_2515# gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X122 vts.t3 vtd.t8 vtd.t9 vts.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X123 vtd.t2 sensor_0.b.t31 gnd.t86 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X124 buffer_0.b buffer_0.b.t9 vd.t34 vd.t33 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X125 out_buff.t3 buffer_0.d gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X126 out_buff.t28 buffer_0.d sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X127 a_16356_5320# a_16190_3988# gnd.t17 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X128 out_buff.t9 buffer_0.d gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X129 vtd.t23 vtd.t22 vts.t1 vts.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X130 vtd.t1 sensor_0.b.t32 gnd.t15 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X131 vd.t82 a_15712_3988# sigma-delta_0.x1.D vd.t81 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X132 sensor_0.c vtd.t27 sensor_0.b.t17 vd.t35 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X133 a_15214_5320# a_15048_3988# gnd.t152 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X134 vd.t84 out.t2 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X135 vd.t32 buffer_0.b.t13 out_buff.t15 vd.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X136 buffer_0.d buffer_0.a.t25 vd.t50 vd.t49 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X137 sensor_0.b.t0 vtd.t28 sensor_0.c vd.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X138 a_17020_5320# a_16854_3988# gnd.t84 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X139 out_buff.t12 buffer_0.b.t14 vd.t26 vd.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X140 gnd.t139 sensor_0.b.t3 sensor_0.b.t4 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X141 sensor_0.d vtd.t29 vd.t46 vd.t45 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X142 buffer_0.d buffer_0.d buffer_0.d gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=2.03 ps=18.1 w=1 l=1
X143 a_14791_2515# a_14625_2515# vpwr.t14 vpwr.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X144 a_14882_5320# a_14716_3988# gnd.t167 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X145 gnd.t171 a_15712_3988# sigma-delta_0.x1.D gnd.t170 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X146 sensor_0.d sensor_0.a.t14 sensor_0.c vd.t79 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X147 buffer_0.a.t3 out_buff.t29 buffer_0.c.t2 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X148 buffer_0.d buffer_0.a.t26 vd.t48 vd.t47 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X149 vts.t20 vts.t17 vts.t19 vts.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X150 ib.t4 ib.t2 ib.t3 gnd.t149 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X151 a_14791_2515# a_14625_2515# gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X152 a_15249_2881# a_14625_2515# a_15141_2515# vpwr.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X153 buffer_0.c.t14 vts.t31 buffer_0.b.t6 gnd.t161 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X154 sensor_0.b.t2 sensor_0.b.t1 gnd.t148 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X155 gnd.t6 sensor_0.b.t33 sensor_0.a.t5 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X156 a_16024_5320# a_15712_3988# gnd.t10 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X157 out_buff.t17 buffer_0.b.t15 vd.t44 vd.t43 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X158 buffer_0.b.t8 vts.t32 buffer_0.c.t13 gnd.t163 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X159 buffer_0.b.t2 vts.t33 buffer_0.c.t12 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X160 vd.t85 out.t1 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X161 vd.t72 buffer_0.b.t16 out_buff.t18 vd.t71 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X162 gnd.t137 out_sigma.t2 out.t0 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X163 vd.t1 buffer_0.b.t17 out_buff.t0 vd.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X164 sensor_0.c sensor_0.a.t15 sensor_0.d vd.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X165 gnd.t151 sensor_0.b.t34 vtd.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X166 out_buff.t20 buffer_0.b.t18 vd.t77 vd.t76 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X167 buffer_0.c.t1 out_buff.t30 buffer_0.a.t7 gnd.t120 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X168 gnd.t38 buffer_0.d buffer_0.d gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X169 gnd.t36 buffer_0.d buffer_0.d gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X170 gnd.t81 a_15881_2489# a_15815_2515# gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X171 out_buff.t1 buffer_0.b.t19 vd.t3 vd.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X172 a_15403_2515# a_15359_2757# a_15237_2515# gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X173 buffer_0.d buffer_0.d gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X174 a_15249_2881# vpwr.t3 vpwr.t5 vpwr.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X175 buffer_0.b.t0 vts.t34 buffer_0.c.t11 gnd.t73 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X176 a_15881_2489# vpwr.t0 vpwr.t2 vpwr.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X177 a_14550_5320# out_buff.t19 gnd.t158 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X178 gnd.t79 a_15881_2489# a_16445_2515# gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X179 sensor_0.a.t4 sensor_0.b.t35 gnd.t150 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X180 vpwr.t19 a_15881_2489# a_16445_2515# vpwr.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X181 buffer_0.a.t4 out_buff.t31 buffer_0.c.t0 gnd.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X182 buffer_0.d buffer_0.d gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X183 gnd.t96 gnd.t93 gnd.t95 gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X184 a_15712_3988# gnd.t169 sky130_fd_pr__cap_mim_m3_1 l=27.2 w=27.2
R0 out_buff.n7 out_buff.t13 30.2161
R1 out_buff.n4 out_buff.t16 29.2293
R2 out_buff.n5 out_buff.t18 28.5655
R3 out_buff.n5 out_buff.t20 28.5655
R4 out_buff.n6 out_buff.t15 28.5655
R5 out_buff.n6 out_buff.t12 28.5655
R6 out_buff.n2 out_buff.t0 28.5655
R7 out_buff.n2 out_buff.t1 28.5655
R8 out_buff.n1 out_buff.t14 28.5655
R9 out_buff.n1 out_buff.t17 28.5655
R10 out_buff.n20 out_buff.t24 26.8319
R11 out_buff.n21 out_buff.t30 25.9449
R12 out_buff.n26 out_buff.t31 25.7428
R13 out_buff.n27 out_buff.t22 25.5407
R14 out_buff.n22 out_buff.t29 25.3386
R15 out_buff.n23 out_buff.t21 25.1365
R16 out_buff.n20 out_buff.t23 24.9306
R17 out_buff.n28 out_buff.t25 24.696
R18 out_buff.n25 out_buff.t27 24.5271
R19 out_buff.n24 out_buff.t26 24.1037
R20 out_buff.n0 out_buff.t4 17.4005
R21 out_buff.n0 out_buff.t10 17.4005
R22 out_buff.n10 out_buff.t5 17.4005
R23 out_buff.n10 out_buff.t2 17.4005
R24 out_buff.n11 out_buff.t6 17.4005
R25 out_buff.n11 out_buff.t9 17.4005
R26 out_buff.n12 out_buff.t8 17.4005
R27 out_buff.n12 out_buff.t11 17.4005
R28 out_buff.n13 out_buff.t7 17.4005
R29 out_buff.n13 out_buff.t3 17.4005
R30 out_buff.n30 out_buff.t19 9.50808
R31 out_buff.n31 out_buff 5.53175
R32 out_buff.n14 out_buff.n13 2.74907
R33 out_buff.n17 out_buff.n9 2.41728
R34 out_buff.n24 out_buff.n23 2.30343
R35 out_buff.n22 out_buff.n21 2.29903
R36 out_buff.n28 out_buff.n27 2.2903
R37 out_buff.n26 out_buff.n25 2.25283
R38 out_buff.n16 out_buff.n15 2.1255
R39 out_buff.n15 out_buff.n14 2.1255
R40 out_buff.n29 out_buff.n19 1.97968
R41 out_buff.n18 out_buff.n17 1.83383
R42 out_buff.n3 out_buff.n1 1.74765
R43 out_buff.n19 out_buff.t28 1.69869
R44 out_buff out_buff.n29 1.51612
R45 out_buff.n29 out_buff.n28 1.24394
R46 out_buff.n31 out_buff.n30 1.11925
R47 out_buff.n8 out_buff.n7 1.04217
R48 out_buff.n4 out_buff.n3 1.0005
R49 out_buff.n9 out_buff.n4 0.938
R50 out_buff.n25 out_buff.n24 0.680308
R51 out_buff.n23 out_buff.n22 0.678839
R52 out_buff.n27 out_buff.n26 0.678839
R53 out_buff.n8 out_buff.n5 0.664316
R54 out_buff.n3 out_buff.n2 0.664316
R55 out_buff.n9 out_buff.n8 0.646333
R56 out_buff.n21 out_buff.n20 0.63023
R57 out_buff.n7 out_buff.n6 0.610444
R58 out_buff.n18 out_buff.n0 0.582399
R59 out_buff.n15 out_buff.n11 0.582399
R60 out_buff.n14 out_buff.n12 0.582399
R61 out_buff.n16 out_buff.n10 0.579923
R62 out_buff.n17 out_buff.n16 0.333833
R63 out_buff out_buff.n31 0.253
R64 out_buff.n19 out_buff.n18 0.250559
R65 out_buff.n30 out_buff 0.05675
R66 gnd.n267 gnd.n264 10830.2
R67 gnd.n137 gnd.n136 6394.13
R68 gnd.n61 gnd.t158 2974.74
R69 gnd.n140 gnd.n137 1867.45
R70 gnd.n137 gnd.t23 1351.39
R71 gnd.n47 gnd.n46 1273.6
R72 gnd.n58 gnd.n57 1260.8
R73 gnd.n54 gnd.n41 1088.88
R74 gnd.n31 gnd.n30 940.25
R75 gnd gnd.n61 642.758
R76 gnd.n206 gnd.n205 585
R77 gnd.n260 gnd.n259 585
R78 gnd.n262 gnd.n261 585
R79 gnd.n165 gnd.n164 585
R80 gnd.n148 gnd.n147 533.923
R81 gnd.t16 gnd.t10 523.77
R82 gnd.n148 gnd.n3 505.849
R83 gnd.n170 gnd.t18 396.608
R84 gnd.n269 gnd.t5 392.344
R85 gnd.t74 gnd.n207 353.962
R86 gnd.t23 gnd.t84 278.673
R87 gnd.t84 gnd.t91 278.673
R88 gnd.t91 gnd.t162 278.673
R89 gnd.t162 gnd.t8 278.673
R90 gnd.t135 gnd.t17 278.673
R91 gnd.t10 gnd.t135 278.673
R92 gnd.t153 gnd.t16 278.673
R93 gnd.t11 gnd.t153 278.673
R94 gnd.t152 gnd.t11 278.673
R95 gnd.t12 gnd.t152 278.673
R96 gnd.t167 gnd.t12 278.673
R97 gnd.t158 gnd.t9 278.673
R98 gnd.t9 gnd.n4 271.957
R99 gnd.n62 gnd.t145 265.026
R100 gnd.n236 gnd.t3 264.406
R101 gnd.n158 gnd.n148 257.24
R102 gnd.t141 gnd.t26 246.649
R103 gnd.n79 gnd.t142 215.036
R104 gnd.t98 gnd.n169 204.702
R105 gnd.n61 gnd.n60 181.864
R106 gnd.t78 gnd.t82 181.843
R107 gnd.t82 gnd.t20 181.843
R108 gnd.n169 gnd.n168 180.179
R109 gnd.n63 gnd.n62 179.542
R110 gnd.n238 gnd.n235 163.766
R111 gnd.t30 gnd.t134 160.564
R112 gnd.n271 gnd.n260 156.236
R113 gnd.n89 gnd.t83 154.317
R114 gnd.n217 gnd.n216 153.976
R115 gnd.n214 gnd.t1 151.393
R116 gnd.t94 gnd.n268 151.393
R117 gnd.n215 gnd.n210 150.648
R118 gnd.n69 gnd.n65 149.835
R119 gnd.n217 gnd.n206 148.707
R120 gnd.t0 gnd.t52 148.462
R121 gnd.t124 gnd.t50 148.462
R122 gnd.t7 gnd.t60 148.462
R123 gnd.t73 gnd.t31 148.462
R124 gnd.t127 gnd.t70 148.462
R125 gnd.t119 gnd.t68 148.462
R126 gnd.t161 gnd.t35 148.462
R127 gnd.t155 gnd.t48 148.462
R128 gnd.t121 gnd.t62 148.462
R129 gnd.t140 gnd.t37 148.462
R130 gnd.t163 gnd.t33 148.462
R131 gnd.t120 gnd.t46 148.462
R132 gnd.t126 gnd.t42 148.462
R133 gnd.t132 gnd.t58 148.462
R134 gnd.t156 gnd.t80 144.12
R135 gnd.n236 gnd.t76 140.732
R136 gnd.t128 gnd.n38 134.233
R137 gnd.n268 gnd.n267 131.137
R138 gnd.n91 gnd.n90 128.757
R139 gnd.t21 gnd.t129 127.677
R140 gnd.n87 gnd.n86 116.754
R141 gnd.n118 gnd.n77 107.24
R142 gnd.n105 gnd.n83 107.24
R143 gnd.t29 gnd.t133 105.43
R144 gnd.n55 gnd.t44 103.922
R145 gnd.t56 gnd.n49 102.686
R146 gnd.t143 gnd.t132 101.448
R147 gnd.t159 gnd.t131 101.448
R148 gnd.n86 gnd.t157 100.001
R149 gnd.n70 gnd.n69 98.6358
R150 gnd.t133 gnd.t21 95.7578
R151 gnd.t145 gnd.t78 93.8233
R152 gnd.n208 gnd.t74 93.8217
R153 gnd.t80 gnd.t29 92.8561
R154 gnd.t134 gnd.t28 92.8561
R155 gnd.t28 gnd.t141 91.8888
R156 gnd.n52 gnd.t40 89.0768
R157 gnd.n35 gnd.n34 88.4582
R158 gnd.n57 gnd.n54 88.0946
R159 gnd.t20 gnd.t156 88.0198
R160 gnd.n44 gnd.t54 85.9839
R161 gnd.n39 gnd.t149 81.6538
R162 gnd.t26 gnd.t24 81.2491
R163 gnd.t5 gnd.n263 76.7633
R164 gnd.n44 gnd.t39 73.6122
R165 gnd.n83 gnd.t130 72.8576
R166 gnd.n86 gnd.t81 70.0005
R167 gnd.t129 gnd.t30 69.6422
R168 gnd.n172 gnd.n165 65.8829
R169 gnd.t24 gnd 62.8715
R170 gnd.n83 gnd.t22 60.5809
R171 gnd.n41 gnd.n37 60.3613
R172 gnd.n52 gnd.t123 59.3847
R173 gnd.t131 gnd.t143 58.1476
R174 gnd.t125 gnd.t159 58.1476
R175 gnd.n90 gnd.t79 57.1434
R176 gnd.n34 gnd.n31 49.4874
R177 gnd.n271 gnd.n262 48.5652
R178 gnd.n49 gnd.t13 45.7758
R179 gnd.n77 gnd.t27 38.5719
R180 gnd.n77 gnd.t25 38.5719
R181 gnd.n252 gnd.t93 37.3602
R182 gnd.n255 gnd.t116 37.3602
R183 gnd.n258 gnd.t101 37.3602
R184 gnd.n177 gnd.t110 37.3602
R185 gnd.n180 gnd.t104 37.3602
R186 gnd.n183 gnd.t113 37.3602
R187 gnd.n107 gnd.n106 34.6358
R188 gnd.n107 gnd.n81 34.6358
R189 gnd.n111 gnd.n81 34.6358
R190 gnd.n112 gnd.n111 34.6358
R191 gnd.n113 gnd.n112 34.6358
R192 gnd.n99 gnd.n98 34.6358
R193 gnd.n100 gnd.n99 34.6358
R194 gnd.n100 gnd.n84 34.6358
R195 gnd.n104 gnd.n84 34.6358
R196 gnd.n94 gnd.n93 34.6358
R197 gnd.n95 gnd.n94 34.6358
R198 gnd.n117 gnd.n79 29.7417
R199 gnd.n93 gnd.n89 27.8593
R200 gnd.n214 gnd.n211 27.7204
R201 gnd.n90 gnd.t146 25.4291
R202 gnd.n158 gnd.t136 25.1825
R203 gnd.n155 gnd.n152 24.9897
R204 gnd.n119 gnd.n118 24.4919
R205 gnd.t168 gnd.n140 23.5887
R206 gnd.n147 gnd.t168 23.5887
R207 gnd.n118 gnd.n117 22.9652
R208 gnd.n39 gnd.t125 19.7952
R209 gnd.n174 gnd.t97 18.6812
R210 gnd.n249 gnd.t107 18.6809
R211 gnd.n95 gnd.n87 17.6946
R212 gnd.n232 gnd.t90 17.4089
R213 gnd.n202 gnd.t139 17.4089
R214 gnd.n243 gnd.t14 17.4084
R215 gnd.n241 gnd.t6 17.4084
R216 gnd.n240 gnd.t85 17.4084
R217 gnd.n243 gnd.t89 17.4084
R218 gnd.n241 gnd.t166 17.4084
R219 gnd.n240 gnd.t150 17.4084
R220 gnd.n232 gnd.t15 17.4079
R221 gnd.n202 gnd.t148 17.4079
R222 gnd.n245 gnd.t77 17.4074
R223 gnd.n245 gnd.t88 17.4074
R224 gnd.n219 gnd.t4 17.4069
R225 gnd.n219 gnd.t2 17.4055
R226 gnd.n248 gnd.t109 17.405
R227 gnd.n248 gnd.t108 17.405
R228 gnd.n251 gnd.t96 17.405
R229 gnd.n251 gnd.t95 17.405
R230 gnd.n254 gnd.t118 17.405
R231 gnd.n254 gnd.t117 17.405
R232 gnd.n257 gnd.t103 17.405
R233 gnd.n257 gnd.t102 17.405
R234 gnd.n173 gnd.t100 17.405
R235 gnd.n173 gnd.t99 17.405
R236 gnd.n176 gnd.t112 17.405
R237 gnd.n176 gnd.t111 17.405
R238 gnd.n179 gnd.t106 17.405
R239 gnd.n179 gnd.t105 17.405
R240 gnd.n182 gnd.t115 17.405
R241 gnd.n182 gnd.t114 17.405
R242 gnd.n73 gnd.t171 17.405
R243 gnd.n221 gnd.t86 17.4034
R244 gnd.n220 gnd.t154 17.4034
R245 gnd.n227 gnd.t92 17.4034
R246 gnd.n226 gnd.t151 17.4034
R247 gnd.n197 gnd.t19 17.4034
R248 gnd.n196 gnd.t75 17.4034
R249 gnd.n191 gnd.t147 17.4034
R250 gnd.n190 gnd.t138 17.4034
R251 gnd.n186 gnd.t72 17.4034
R252 gnd.n185 gnd.t165 17.4034
R253 gnd.n24 gnd.t144 17.4005
R254 gnd.n24 gnd.t160 17.4005
R255 gnd.n22 gnd.t43 17.4005
R256 gnd.n22 gnd.t59 17.4005
R257 gnd.n20 gnd.t34 17.4005
R258 gnd.n20 gnd.t47 17.4005
R259 gnd.n18 gnd.t63 17.4005
R260 gnd.n18 gnd.t38 17.4005
R261 gnd.n16 gnd.t67 17.4005
R262 gnd.n16 gnd.t65 17.4005
R263 gnd.n14 gnd.t41 17.4005
R264 gnd.n14 gnd.t57 17.4005
R265 gnd.n12 gnd.t49 17.4005
R266 gnd.n12 gnd.t45 17.4005
R267 gnd.n10 gnd.t69 17.4005
R268 gnd.n10 gnd.t36 17.4005
R269 gnd.n8 gnd.t32 17.4005
R270 gnd.n8 gnd.t71 17.4005
R271 gnd.n6 gnd.t51 17.4005
R272 gnd.n6 gnd.t61 17.4005
R273 gnd.n5 gnd.t55 17.4005
R274 gnd.n5 gnd.t53 17.4005
R275 gnd.n113 gnd.n79 14.6829
R276 gnd.n38 gnd.t64 14.228
R277 gnd.n269 gnd.t94 12.7943
R278 gnd.t50 gnd.t0 11.135
R279 gnd.t60 gnd.t124 11.135
R280 gnd.t31 gnd.t7 11.135
R281 gnd.t70 gnd.t73 11.135
R282 gnd.t68 gnd.t127 11.135
R283 gnd.t35 gnd.t119 11.135
R284 gnd.t48 gnd.t161 11.135
R285 gnd.t44 gnd.t155 11.135
R286 gnd.t40 gnd.t122 11.135
R287 gnd.t123 gnd.t56 11.135
R288 gnd.t13 gnd.t66 11.135
R289 gnd.t64 gnd.t87 11.135
R290 gnd.t62 gnd.t128 11.135
R291 gnd.t37 gnd.t121 11.135
R292 gnd.t33 gnd.t140 11.135
R293 gnd.t46 gnd.t163 11.135
R294 gnd.t42 gnd.t120 11.135
R295 gnd.t58 gnd.t126 11.135
R296 gnd.n91 gnd.n89 10.9075
R297 gnd.n73 gnd.n72 9.33321
R298 gnd.n172 gnd.n171 9.3005
R299 gnd.n171 gnd.n170 9.3005
R300 gnd.n217 gnd.n209 9.3005
R301 gnd.n209 gnd.n208 9.3005
R302 gnd.n238 gnd.n237 9.3005
R303 gnd.n237 gnd.n236 9.3005
R304 gnd.n271 gnd.n270 9.3005
R305 gnd.n270 gnd.n269 9.3005
R306 gnd.n162 gnd.t137 8.70236
R307 gnd.n170 gnd.t98 8.5297
R308 gnd.n106 gnd.n105 7.90638
R309 gnd.n4 gnd.t167 6.71549
R310 gnd.n35 gnd.t164 4.94919
R311 gnd.n115 gnd.n79 4.6505
R312 gnd.n93 gnd.n92 4.6505
R313 gnd.n94 gnd.n88 4.6505
R314 gnd.n96 gnd.n95 4.6505
R315 gnd.n98 gnd.n97 4.6505
R316 gnd.n99 gnd.n85 4.6505
R317 gnd.n101 gnd.n100 4.6505
R318 gnd.n102 gnd.n84 4.6505
R319 gnd.n104 gnd.n103 4.6505
R320 gnd.n106 gnd.n82 4.6505
R321 gnd.n108 gnd.n107 4.6505
R322 gnd.n109 gnd.n81 4.6505
R323 gnd.n111 gnd.n110 4.6505
R324 gnd.n112 gnd.n80 4.6505
R325 gnd.n114 gnd.n113 4.6505
R326 gnd.n117 gnd.n116 4.6505
R327 gnd.n118 gnd.n78 4.6505
R328 gnd.n75 gnd.n74 4.5005
R329 gnd.n76 gnd.n74 4.5005
R330 gnd gnd.n122 3.79922
R331 gnd.n123 gnd.n0 3.24248
R332 gnd.n26 gnd.n0 3.01925
R333 gnd.n126 gnd.n124 2.6505
R334 gnd.n98 gnd.n87 2.63579
R335 gnd gnd.n162 2.5773
R336 gnd.n120 gnd.n74 2.25328
R337 gnd.n105 gnd.n104 1.88285
R338 gnd.n163 gnd 1.8224
R339 gnd.n7 gnd.n5 1.66573
R340 gnd.n124 gnd.t169 1.47915
R341 gnd.n25 gnd.n23 1.3755
R342 gnd.n163 gnd.n0 1.30732
R343 gnd.n124 gnd.n123 1.22706
R344 gnd.n9 gnd.n7 1.08383
R345 gnd.n13 gnd.n11 1.08383
R346 gnd.n15 gnd.n13 1.08383
R347 gnd.n17 gnd.n15 1.08383
R348 gnd.n21 gnd.n19 1.08383
R349 gnd.n23 gnd.n21 1.08383
R350 gnd.n11 gnd.n9 1.04217
R351 gnd.n19 gnd.n17 1.04217
R352 gnd.n23 gnd.n22 0.582399
R353 gnd.n21 gnd.n20 0.582399
R354 gnd.n19 gnd.n18 0.582399
R355 gnd.n17 gnd.n16 0.582399
R356 gnd.n15 gnd.n14 0.582399
R357 gnd.n13 gnd.n12 0.582399
R358 gnd.n11 gnd.n10 0.582399
R359 gnd.n7 gnd.n6 0.582399
R360 gnd.n9 gnd.n8 0.579923
R361 gnd.n25 gnd.n24 0.57713
R362 gnd.n130 gnd.n71 0.54125
R363 gnd.n71 gnd.n70 0.541165
R364 gnd.n225 gnd.n219 0.447415
R365 gnd.n231 gnd.n225 0.438
R366 gnd.n233 gnd.n231 0.438
R367 gnd.n275 gnd.n274 0.401236
R368 gnd.n27 gnd.n25 0.392443
R369 gnd.n195 gnd.n189 0.375501
R370 gnd.n234 gnd.n233 0.375501
R371 gnd.n201 gnd.n195 0.3755
R372 gnd.n203 gnd.n201 0.3755
R373 gnd.n242 gnd.n240 0.373217
R374 gnd.n244 gnd.n242 0.371401
R375 gnd.n246 gnd.n244 0.369555
R376 gnd.n159 gnd.n2 0.366293
R377 gnd.n150 gnd.n149 0.365897
R378 gnd.n158 gnd.n150 0.365897
R379 gnd.n2 gnd.n1 0.365897
R380 gnd.n135 gnd.n134 0.347558
R381 gnd.n134 gnd.n133 0.347269
R382 gnd.n247 gnd.n246 0.338503
R383 gnd.n204 gnd.n203 0.330858
R384 gnd.n204 gnd.n184 0.290469
R385 gnd.n37 gnd.n36 0.288252
R386 gnd.n36 gnd.n35 0.288252
R387 gnd.n234 gnd.n218 0.281539
R388 gnd.n27 gnd.n26 0.274914
R389 gnd.n239 gnd.n234 0.245825
R390 gnd.n273 gnd.n247 0.244548
R391 gnd.n275 gnd.n163 0.230614
R392 gnd.n247 gnd.n239 0.180349
R393 gnd.n218 gnd.n204 0.156539
R394 gnd.n92 gnd.n91 0.144332
R395 gnd.n142 gnd.n141 0.1305
R396 gnd.t168 gnd.n142 0.1305
R397 gnd.n144 gnd.n143 0.1305
R398 gnd.t168 gnd.n144 0.1305
R399 gnd.n92 gnd.n88 0.120292
R400 gnd.n96 gnd.n88 0.120292
R401 gnd.n97 gnd.n96 0.120292
R402 gnd.n97 gnd.n85 0.120292
R403 gnd.n101 gnd.n85 0.120292
R404 gnd.n102 gnd.n101 0.120292
R405 gnd.n103 gnd.n102 0.120292
R406 gnd.n103 gnd.n82 0.120292
R407 gnd.n108 gnd.n82 0.120292
R408 gnd.n109 gnd.n108 0.120292
R409 gnd.n110 gnd.n109 0.120292
R410 gnd.n110 gnd.n80 0.120292
R411 gnd.n114 gnd.n80 0.120292
R412 gnd.n115 gnd.n114 0.120292
R413 gnd.n116 gnd.n115 0.120292
R414 gnd.n116 gnd.n78 0.120292
R415 gnd.n154 gnd.n153 0.10956
R416 gnd.n157 gnd.n156 0.10956
R417 gnd.t136 gnd.n157 0.10956
R418 gnd.n67 gnd.n66 0.10956
R419 gnd.t170 gnd.n67 0.10956
R420 gnd.n68 gnd.t170 0.10956
R421 gnd.n69 gnd.n68 0.10956
R422 gnd.n155 gnd.n154 0.109112
R423 gnd.n135 gnd.n132 0.0849523
R424 gnd.n132 gnd.n131 0.0845034
R425 gnd.n276 gnd.n275 0.0772045
R426 gnd.n276 gnd 0.0755
R427 gnd.n78 gnd.n75 0.0734167
R428 gnd.n250 gnd.n249 0.073412
R429 gnd.n175 gnd.n174 0.0734113
R430 gnd.n26 gnd 0.06925
R431 gnd.n176 gnd.n175 0.0610469
R432 gnd.n177 gnd.n176 0.0610469
R433 gnd.n179 gnd.n178 0.0610469
R434 gnd.n180 gnd.n179 0.0610469
R435 gnd.n182 gnd.n181 0.0610469
R436 gnd.n183 gnd.n182 0.0610469
R437 gnd.n251 gnd.n250 0.0610469
R438 gnd.n252 gnd.n251 0.0610469
R439 gnd.n254 gnd.n253 0.0610469
R440 gnd.n255 gnd.n254 0.0610469
R441 gnd.n257 gnd.n256 0.0610469
R442 gnd.n258 gnd.n257 0.0610469
R443 gnd.n272 gnd.n258 0.0573558
R444 gnd.n184 gnd.n183 0.0573547
R445 gnd.n273 gnd.n272 0.0464211
R446 gnd.n178 gnd.n177 0.0426875
R447 gnd.n181 gnd.n180 0.0426875
R448 gnd.n253 gnd.n252 0.0426875
R449 gnd.n256 gnd.n255 0.0426875
R450 gnd.n65 gnd.n64 0.0425017
R451 gnd.n64 gnd.n63 0.0425017
R452 gnd.n29 gnd.n28 0.0425017
R453 gnd.n31 gnd.n29 0.0425017
R454 gnd.n46 gnd.n45 0.0425017
R455 gnd.n45 gnd.n44 0.0425017
R456 gnd.n33 gnd.n32 0.0425017
R457 gnd.n34 gnd.n33 0.0425017
R458 gnd.n59 gnd.n58 0.0425017
R459 gnd.n60 gnd.n59 0.0425017
R460 gnd.n274 gnd 0.0395625
R461 gnd gnd.n276 0.0345909
R462 gnd.n76 gnd 0.0330521
R463 gnd.n123 gnd 0.03175
R464 gnd.n174 gnd.n173 0.031274
R465 gnd.n249 gnd.n248 0.0312734
R466 gnd.n121 gnd.n75 0.0265417
R467 gnd.n152 gnd.n151 0.0264102
R468 gnd.n119 gnd 0.0226354
R469 gnd.n233 gnd.n232 0.0153409
R470 gnd.n230 gnd.n228 0.0129048
R471 gnd.n121 gnd.n120 0.0114272
R472 gnd.n224 gnd.n222 0.0114167
R473 gnd.n120 gnd.n119 0.0113582
R474 gnd.n122 gnd.n74 0.0110001
R475 gnd.n216 gnd.n215 0.0092427
R476 gnd.n215 gnd.n214 0.0092427
R477 gnd.n266 gnd.n265 0.00883856
R478 gnd.n267 gnd.n266 0.00883856
R479 gnd.n167 gnd.n166 0.00883856
R480 gnd.n168 gnd.n167 0.00883856
R481 gnd.n127 gnd.n73 0.00867757
R482 gnd.n203 gnd.n202 0.00792873
R483 gnd.n146 gnd.n145 0.00762598
R484 gnd.n147 gnd.n146 0.00762598
R485 gnd.n139 gnd.n138 0.00762598
R486 gnd.n140 gnd.n139 0.00762598
R487 gnd.n127 gnd.n126 0.00634112
R488 gnd gnd.n76 0.00570833
R489 gnd.n200 gnd.n198 0.00546432
R490 gnd.n187 gnd.n185 0.00502806
R491 gnd.n192 gnd.n190 0.00502806
R492 gnd.n198 gnd.n196 0.00502805
R493 gnd.n222 gnd.n220 0.00502803
R494 gnd.n228 gnd.n226 0.00502803
R495 gnd.n57 gnd.n56 0.00498892
R496 gnd.n56 gnd.n55 0.00498892
R497 gnd.n213 gnd.n212 0.00487141
R498 gnd.n214 gnd.n213 0.00487141
R499 gnd.n54 gnd.n53 0.00466542
R500 gnd.n53 gnd.n52 0.00466542
R501 gnd.n130 gnd.n129 0.00441022
R502 gnd.n187 gnd.n186 0.00402807
R503 gnd.n192 gnd.n191 0.00402806
R504 gnd.n198 gnd.n197 0.00402806
R505 gnd.n222 gnd.n221 0.00402804
R506 gnd.n228 gnd.n227 0.00402803
R507 gnd.n194 gnd.n192 0.00397623
R508 gnd.n129 gnd.n128 0.00391284
R509 gnd.n128 gnd.n127 0.00391159
R510 gnd.n43 gnd.n42 0.00271942
R511 gnd.n49 gnd.n43 0.00271942
R512 gnd.n48 gnd.n47 0.00271942
R513 gnd.n49 gnd.n48 0.00271942
R514 gnd.n51 gnd.n50 0.00258271
R515 gnd.n52 gnd.n51 0.00258271
R516 gnd.n189 gnd.n187 0.00248813
R517 gnd.n274 gnd.n273 0.00245312
R518 gnd.n160 gnd.n159 0.00236777
R519 gnd.t136 gnd.n155 0.00194448
R520 gnd.n41 gnd.n40 0.00190526
R521 gnd.n40 gnd.n39 0.00190526
R522 gnd.n161 gnd.n160 0.00186816
R523 gnd.n272 gnd.n271 0.00152216
R524 gnd.n184 gnd.n172 0.00152195
R525 gnd.n230 gnd.n229 0.00138337
R526 gnd.n224 gnd.n223 0.00138109
R527 gnd.n200 gnd.n199 0.00134613
R528 gnd.n194 gnd.n193 0.00134049
R529 gnd.n189 gnd.n188 0.001335
R530 gnd.n162 gnd.n161 0.00124275
R531 gnd.n244 gnd.n243 0.00121065
R532 gnd.n242 gnd.n241 0.001204
R533 gnd.n136 gnd.n135 0.00104118
R534 gnd.n122 gnd.n121 0.00100955
R535 gnd.n136 gnd.n130 0.00100261
R536 gnd.n246 gnd.n245 0.00100079
R537 gnd.n159 gnd.n158 0.00100039
R538 gnd.n218 gnd.n217 0.000522345
R539 gnd.n239 gnd.n238 0.000522345
R540 gnd.n126 gnd.n125 0.00051897
R541 gnd.n41 gnd.n27 0.000503131
R542 gnd.n231 gnd.n230 0.000501021
R543 gnd.n225 gnd.n224 0.000501021
R544 gnd.n195 gnd.n194 0.000500672
R545 gnd.n201 gnd.n200 0.000500672
R546 buffer_0.a.n6 buffer_0.a.t26 40.2461
R547 buffer_0.a.n2 buffer_0.a.t21 40.2461
R548 buffer_0.a.n10 buffer_0.a.t10 39.5292
R549 buffer_0.a.n9 buffer_0.a.t20 39.5292
R550 buffer_0.a.n8 buffer_0.a.t17 39.5292
R551 buffer_0.a.n7 buffer_0.a.t25 39.5292
R552 buffer_0.a.n6 buffer_0.a.t18 39.5292
R553 buffer_0.a.n5 buffer_0.a.t19 39.5292
R554 buffer_0.a.n4 buffer_0.a.t24 39.5292
R555 buffer_0.a.n3 buffer_0.a.t23 39.5292
R556 buffer_0.a.n2 buffer_0.a.t22 39.5292
R557 buffer_0.a.n12 buffer_0.a.t11 28.576
R558 buffer_0.a.n1 buffer_0.a.t14 25.2845
R559 buffer_0.a.n0 buffer_0.a.t12 24.699
R560 buffer_0.a.n1 buffer_0.a.t16 17.4081
R561 buffer_0.a.n1 buffer_0.a.t1 17.4005
R562 buffer_0.a.n1 buffer_0.a.t15 17.4005
R563 buffer_0.a.n17 buffer_0.a.t9 17.4005
R564 buffer_0.a.n17 buffer_0.a.t3 17.4005
R565 buffer_0.a.n15 buffer_0.a.t0 17.4005
R566 buffer_0.a.n15 buffer_0.a.t6 17.4005
R567 buffer_0.a.n13 buffer_0.a.t8 17.4005
R568 buffer_0.a.n13 buffer_0.a.t4 17.4005
R569 buffer_0.a.n0 buffer_0.a.t13 17.4005
R570 buffer_0.a.n0 buffer_0.a.t5 17.4005
R571 buffer_0.a.n19 buffer_0.a.t7 17.4005
R572 buffer_0.a.n19 buffer_0.a.t2 17.4005
R573 buffer_0.a.n14 buffer_0.a.n0 2.76905
R574 buffer_0.a.n20 buffer_0.a.n1 2.69153
R575 buffer_0.a.n16 buffer_0.a.n14 2.16717
R576 buffer_0.a.n18 buffer_0.a.n16 2.1255
R577 buffer_0.a.n21 buffer_0.a.n20 1.2505
R578 buffer_0.a.n10 buffer_0.a.n9 1.06739
R579 buffer_0.a.n21 buffer_0.a.n18 0.917167
R580 buffer_0.a buffer_0.a.n12 0.862147
R581 buffer_0.a.n11 buffer_0.a.n5 0.749569
R582 buffer_0.a.n7 buffer_0.a.n6 0.717388
R583 buffer_0.a.n8 buffer_0.a.n7 0.717388
R584 buffer_0.a.n9 buffer_0.a.n8 0.717388
R585 buffer_0.a.n3 buffer_0.a.n2 0.717388
R586 buffer_0.a.n4 buffer_0.a.n3 0.717388
R587 buffer_0.a.n5 buffer_0.a.n4 0.717388
R588 buffer_0.a.n20 buffer_0.a.n19 0.526026
R589 buffer_0.a.n16 buffer_0.a.n15 0.52595
R590 buffer_0.a buffer_0.a.n21 0.521392
R591 buffer_0.a.n18 buffer_0.a.n17 0.516495
R592 buffer_0.a.n14 buffer_0.a.n13 0.516495
R593 buffer_0.a.n11 buffer_0.a.n10 0.349569
R594 buffer_0.a.n12 buffer_0.a.n11 0.271856
R595 vd.n62 vd.n59 2142.35
R596 vd.n31 vd.n28 1304.47
R597 vd.n66 vd.n60 1164.71
R598 vd.n68 vd.n56 1164.71
R599 vd.n44 vd.n36 1070.68
R600 vd.n68 vd.n57 977.648
R601 vd.n66 vd.n59 952.942
R602 vd.t71 vd.t33 537.318
R603 vd.t33 vd.t37 526.24
R604 vd.t61 vd.t63 526.24
R605 vd.t59 vd.t61 512.391
R606 vd.t22 vd.t29 357.289
R607 vd.t29 vd.t43 357.289
R608 vd.t43 vd.t0 357.289
R609 vd.t37 vd.t2 357.289
R610 vd.t76 vd.t71 357.289
R611 vd.t31 vd.t76 357.289
R612 vd.t25 vd.t31 357.289
R613 vd.t57 vd.t55 357.289
R614 vd.t55 vd.t53 357.289
R615 vd.t53 vd.t51 357.289
R616 vd.t67 vd.t59 357.289
R617 vd.t49 vd.t67 357.289
R618 vd.t65 vd.t49 357.289
R619 vd.n27 vd.t22 354.529
R620 vd.n34 vd.t57 282.507
R621 vd.n34 vd.t27 254.811
R622 vd.n64 vd.n63 228.518
R623 vd.n63 vd.n54 228.518
R624 vd.n43 vd.n40 223.625
R625 vd.n128 vd.n125 206.306
R626 vd.n37 vd.t47 204.957
R627 vd.n96 vd.n95 168.66
R628 vd.t6 vd.n109 156.245
R629 vd.n37 vd.t65 152.333
R630 vd.n67 vd.t81 144.606
R631 vd.n29 vd.t25 144.024
R632 vd.n91 vd.t35 143.697
R633 vd.n113 vd.t73 143.697
R634 vd.n135 vd.n132 142.306
R635 vd.n62 vd.n61 135.465
R636 vd.n36 vd.n31 127.248
R637 vd.n115 vd.n112 126.871
R638 vd.n44 vd.n43 117.835
R639 vd.n88 vd.n87 111.421
R640 vd.n69 vd.n54 104.282
R641 vd.n65 vd.n64 101.647
R642 vd.n41 vd.t14 92.7848
R643 vd.n133 vd.t36 86.6752
R644 vd.n96 vd.n90 85.0829
R645 vd.n126 vd.t10 71.8492
R646 vd.n91 vd.t18 65.0065
R647 vd.n84 vd.t17 63.6934
R648 vd.n98 vd.t9 63.6821
R649 vd.n104 vd.t5 63.6292
R650 vd.n128 vd.n122 63.2476
R651 vd.n133 vd.t39 60.4447
R652 vd.t36 vd.t69 58.1638
R653 vd.t10 vd.t75 58.1638
R654 vd.n120 vd.t45 42.1974
R655 vd.n123 vd.t78 42.1974
R656 vd.n70 vd.n69 31.105
R657 vd.n20 vd.t62 29.2512
R658 vd.n15 vd.t58 29.2303
R659 vd.n10 vd.t72 29.2303
R660 vd.n9 vd.t34 29.2303
R661 vd.n26 vd.t16 28.5795
R662 vd.n3 vd.t30 28.57
R663 vd.n23 vd.t50 28.5655
R664 vd.n23 vd.t66 28.5655
R665 vd.n21 vd.t60 28.5655
R666 vd.n21 vd.t68 28.5655
R667 vd.n18 vd.t52 28.5655
R668 vd.n18 vd.t64 28.5655
R669 vd.n16 vd.t56 28.5655
R670 vd.n16 vd.t54 28.5655
R671 vd.n13 vd.t26 28.5655
R672 vd.n13 vd.t28 28.5655
R673 vd.n11 vd.t77 28.5655
R674 vd.n11 vd.t32 28.5655
R675 vd.n7 vd.t3 28.5655
R676 vd.n7 vd.t38 28.5655
R677 vd.n5 vd.t44 28.5655
R678 vd.n5 vd.t1 28.5655
R679 vd.n25 vd.t48 28.5655
R680 vd.n25 vd.t15 28.5655
R681 vd.n93 vd.t4 28.5119
R682 vd.n65 vd.n48 27.9188
R683 vd.n106 vd.n101 24.5501
R684 vd.n70 vd.n53 22.401
R685 vd.n78 vd.n77 22.4005
R686 vd.n53 vd.n51 22.4005
R687 vd.n110 vd.t6 21.0989
R688 vd.n4 vd.t21 19.8115
R689 vd.n26 vd.t13 19.8115
R690 vd.t45 vd.t24 19.3883
R691 vd.n79 vd.n48 19.201
R692 vd.n79 vd.n78 19.2005
R693 vd.n126 vd.t79 17.1073
R694 vd.n97 vd.t46 14.5056
R695 vd.n83 vd.t70 14.472
R696 vd.n97 vd.t11 14.4415
R697 vd.n99 vd.t12 14.4153
R698 vd.n85 vd.t19 14.4127
R699 vd.n103 vd.t7 14.4041
R700 vd.n83 vd.t20 14.3878
R701 vd.n101 vd.t8 14.2867
R702 vd.n3 vd.t23 14.2847
R703 vd.n102 vd.t74 14.283
R704 vd.n102 vd.t41 14.283
R705 vd.t18 vd.t42 11.4051
R706 vd.n55 vd.n51 10.5605
R707 vd.n77 vd.n50 9.6005
R708 vd.n2 vd.t80 9.5742
R709 vd.n74 vd.t82 9.52337
R710 vd.n106 vd.n105 9.3005
R711 vd.n107 vd.n106 4.5005
R712 vd.n141 vd.n140 3.73002
R713 vd.n113 vd.t40 3.42187
R714 vd vd.n82 2.438
R715 vd.n55 vd.n50 2.2405
R716 vd.n139 vd 2.08242
R717 vd vd.n107 1.83279
R718 vd.n6 vd.n4 1.47391
R719 vd vd.n26 1.0363
R720 vd.n9 vd.n8 1.0005
R721 vd.n20 vd.n19 1.0005
R722 vd.n138 vd.n85 0.862412
R723 vd.n139 vd.n138 0.834744
R724 vd.n8 vd.n6 0.813
R725 vd.n12 vd.n10 0.813
R726 vd.n19 vd.n17 0.813
R727 vd.n14 vd.n12 0.78175
R728 vd.n17 vd.n15 0.78175
R729 vd.n24 vd.n22 0.78175
R730 vd.n103 vd.n102 0.721906
R731 vd.n24 vd.n23 0.665316
R732 vd.n22 vd.n21 0.665316
R733 vd.n19 vd.n18 0.665316
R734 vd.n14 vd.n13 0.665316
R735 vd.n12 vd.n11 0.665316
R736 vd.n8 vd.n7 0.665316
R737 vd.n6 vd.n5 0.665316
R738 vd.n15 vd.n14 0.6255
R739 vd.n17 vd.n16 0.611443
R740 vd.n104 vd.n103 0.608294
R741 vd.n22 vd.n20 0.59425
R742 vd.n117 vd.n99 0.576317
R743 vd.n137 vd.n136 0.5755
R744 vd.n136 vd.n129 0.488
R745 vd.n117 vd.n116 0.463
R746 vd.n99 vd.n98 0.344245
R747 vd.n46 vd.n24 0.302583
R748 vd.n116 vd 0.2755
R749 vd.n129 vd.n117 0.238
R750 vd.n140 vd.n46 0.23013
R751 vd.n10 vd.n9 0.21925
R752 vd.n142 vd.n141 0.2005
R753 vd.n72 vd.n71 0.146341
R754 vd.n72 vd.n47 0.146333
R755 vd.n66 vd.n65 0.130052
R756 vd.n67 vd.n66 0.130052
R757 vd.n84 vd.n83 0.129979
R758 vd.n82 vd.n47 0.1255
R759 vd.n142 vd 0.1255
R760 vd.n101 vd.n100 0.122252
R761 vd.n105 vd.n104 0.116172
R762 vd.n69 vd.n68 0.107375
R763 vd.n68 vd.n67 0.107375
R764 vd.n142 vd.n2 0.0822638
R765 vd.n0 vd.t83 0.0686501
R766 vd.n1 vd.n0 0.06865
R767 vd.n140 vd.n139 0.0648158
R768 vd.n76 vd.n49 0.0456031
R769 vd.n73 vd.n52 0.0456031
R770 vd.n71 vd.n52 0.0456031
R771 vd.n45 vd 0.0421667
R772 vd.n81 vd.n80 0.0391598
R773 vd.n80 vd.n49 0.0391598
R774 vd.n141 vd 0.0372647
R775 vd.n64 vd.n59 0.0349892
R776 vd.n59 vd.t81 0.0349892
R777 vd.n57 vd.n54 0.0349892
R778 vd.n61 vd.n57 0.0333079
R779 vd.n98 vd.n97 0.0321654
R780 vd.n90 vd.n89 0.0307238
R781 vd.n89 vd.n88 0.0302348
R782 vd.n85 vd.n84 0.0267443
R783 vd.n74 vd.n73 0.0217629
R784 vd.n76 vd.n75 0.0198299
R785 vd.n107 vd.n100 0.0176875
R786 vd.n112 vd.n111 0.0175052
R787 vd.n111 vd.n110 0.0175052
R788 vd.n43 vd.n42 0.0168558
R789 vd.n42 vd.n41 0.0168558
R790 vd.n132 vd.n131 0.0150968
R791 vd.n131 vd.n130 0.0150968
R792 vd vd.n142 0.013
R793 vd.n58 vd.n56 0.0125538
R794 vd.n95 vd.n94 0.0122827
R795 vd.n94 vd.n93 0.0122827
R796 vd.n56 vd.n55 0.0120596
R797 vd.n46 vd.n45 0.0109167
R798 vd.n105 vd.n100 0.009875
R799 vd.n40 vd.n39 0.00979742
R800 vd.n28 vd.n27 0.00979742
R801 vd.n125 vd.n124 0.00973799
R802 vd.n124 vd.n123 0.00973799
R803 vd.n2 vd.n1 0.00846782
R804 vd.n138 vd.n137 0.00675
R805 vd.n63 vd.n62 0.00627981
R806 vd.n44 vd.n38 0.0055
R807 vd.n38 vd.n37 0.0055
R808 vd.n75 vd.n74 0.00501031
R809 vd.n4 vd.n3 0.00500317
R810 vd.n26 vd.n25 0.00454578
R811 vd.n135 vd.n134 0.00391284
R812 vd.n134 vd.n133 0.00391284
R813 vd.n128 vd.n127 0.00391284
R814 vd.n127 vd.n126 0.00391284
R815 vd.n115 vd.n114 0.00391284
R816 vd.n114 vd.n113 0.00391284
R817 vd.n96 vd.n92 0.00391284
R818 vd.n92 vd.n91 0.00391284
R819 vd.n109 vd.n108 0.00347027
R820 vd.n87 vd.n86 0.00347027
R821 vd.n61 vd.t81 0.00318081
R822 vd.n122 vd.n121 0.00275116
R823 vd.n121 vd.n120 0.00275116
R824 vd.n31 vd.n30 0.00186586
R825 vd.n30 vd.n29 0.00186586
R826 vd.n60 vd.n58 0.0018171
R827 vd.n36 vd.n35 0.00173262
R828 vd.n35 vd.n34 0.00173262
R829 vd.n120 vd.n119 0.00162558
R830 vd.n119 vd.n118 0.00162558
R831 vd.n60 vd.n50 0.00131751
R832 vd.n75 vd.n50 0.00131744
R833 vd.n80 vd.n79 0.00119114
R834 vd.n33 vd.n32 0.00111631
R835 vd.n34 vd.n33 0.00111631
R836 vd.n81 vd.n48 0.00101609
R837 vd.n67 vd.n58 0.00100038
R838 vd.n71 vd.n70 0.00100009
R839 vd.n53 vd.n52 0.000659706
R840 vd.n77 vd.n76 0.000659706
R841 vd.n78 vd.n49 0.000543686
R842 vd.n73 vd.n51 0.000543686
R843 vd.n136 vd.n135 0.000532663
R844 vd.n129 vd.n128 0.000532663
R845 vd.n116 vd.n115 0.000532663
R846 vd.n137 vd.n96 0.000532663
R847 vd.n45 vd.n44 0.000511142
R848 vd.n82 vd.n81 0.000507883
R849 vd.n49 vd.n47 0.000507883
R850 vd.n73 vd.n72 0.000507883
R851 vd.n0 vd.t85 0.000500086
R852 vd.n1 vd.t84 0.000500086
R853 sensor_0.b.t9 sensor_0.b.t1 74.8549
R854 sensor_0.b.t7 sensor_0.b.t9 74.8549
R855 sensor_0.b.t15 sensor_0.b.t7 74.8549
R856 sensor_0.b.t11 sensor_0.b.t3 74.8549
R857 sensor_0.b.t5 sensor_0.b.t11 74.8549
R858 sensor_0.b.t13 sensor_0.b.t5 74.8549
R859 sensor_0.b.t24 sensor_0.b.t32 74.8549
R860 sensor_0.b.t31 sensor_0.b.t24 74.8549
R861 sensor_0.b.t23 sensor_0.b.t31 74.8549
R862 sensor_0.b.t34 sensor_0.b.t26 74.8549
R863 sensor_0.b.t21 sensor_0.b.t34 74.8549
R864 sensor_0.b.t29 sensor_0.b.t21 74.8549
R865 sensor_0.b.t27 sensor_0.b.t20 74.8549
R866 sensor_0.b.t28 sensor_0.b.t27 74.8549
R867 sensor_0.b.t35 sensor_0.b.t28 74.8549
R868 sensor_0.b.t22 sensor_0.b.t30 74.8549
R869 sensor_0.b.t33 sensor_0.b.t22 74.8549
R870 sensor_0.b.t25 sensor_0.b.t33 74.8549
R871 sensor_0.b.n7 sensor_0.b.t25 38.3763
R872 sensor_0.b.n11 sensor_0.b.t15 37.3627
R873 sensor_0.b.n10 sensor_0.b.t13 37.3602
R874 sensor_0.b.n9 sensor_0.b.t23 37.3602
R875 sensor_0.b.n8 sensor_0.b.t29 37.3602
R876 sensor_0.b.n7 sensor_0.b.t35 37.3602
R877 sensor_0.b.n12 sensor_0.b.t2 18.2715
R878 sensor_0.b.n3 sensor_0.b.t4 18.1717
R879 sensor_0.b.n14 sensor_0.b.t16 17.427
R880 sensor_0.b.n13 sensor_0.b.t8 17.4116
R881 sensor_0.b.n3 sensor_0.b.t12 17.4101
R882 sensor_0.b.n12 sensor_0.b.t10 17.4101
R883 sensor_0.b.n4 sensor_0.b.t6 17.4058
R884 sensor_0.b.n5 sensor_0.b.t14 17.4056
R885 sensor_0.b.n0 sensor_0.b.t17 14.283
R886 sensor_0.b.n0 sensor_0.b.t0 14.283
R887 sensor_0.b.n1 sensor_0.b.t18 14.283
R888 sensor_0.b.n1 sensor_0.b.t19 14.283
R889 sensor_0.b.n6 sensor_0.b.n5 3.22928
R890 sensor_0.b.n6 sensor_0.b.n2 2.2255
R891 sensor_0.b.n11 sensor_0.b.n10 1.01759
R892 sensor_0.b.n8 sensor_0.b.n7 1.01657
R893 sensor_0.b.n9 sensor_0.b.n8 1.01657
R894 sensor_0.b.n10 sensor_0.b.n9 1.01657
R895 sensor_0.b.n13 sensor_0.b.n12 0.865287
R896 sensor_0.b sensor_0.b.n15 0.851048
R897 sensor_0.b.n14 sensor_0.b.n13 0.777059
R898 sensor_0.b.n5 sensor_0.b.n4 0.718555
R899 sensor_0.b.n4 sensor_0.b.n3 0.710921
R900 sensor_0.b.n2 sensor_0.b.n0 0.49917
R901 sensor_0.b sensor_0.b.n6 0.341125
R902 sensor_0.b.n15 sensor_0.b.n14 0.325292
R903 sensor_0.b.n15 sensor_0.b.n11 0.202053
R904 sensor_0.b.n2 sensor_0.b.n1 0.17167
R905 sensor_0.a.n2 sensor_0.a.t15 64.1667
R906 sensor_0.a.n0 sensor_0.a.t0 63.6292
R907 sensor_0.a.n4 sensor_0.a.t13 63.6292
R908 sensor_0.a.n3 sensor_0.a.t12 63.6292
R909 sensor_0.a.n2 sensor_0.a.t14 63.6292
R910 sensor_0.a.n1 sensor_0.a.t2 63.6275
R911 sensor_0.a.n8 sensor_0.a.t6 18.2715
R912 sensor_0.a.n5 sensor_0.a.t11 18.2714
R913 sensor_0.a.n10 sensor_0.a.t9 17.4132
R914 sensor_0.a.n7 sensor_0.a.t4 17.4132
R915 sensor_0.a.n6 sensor_0.a.t7 17.4116
R916 sensor_0.a.n8 sensor_0.a.t10 17.4101
R917 sensor_0.a.n5 sensor_0.a.t8 17.4101
R918 sensor_0.a.n9 sensor_0.a.t5 17.4057
R919 sensor_0.a.n1 sensor_0.a.t3 14.5343
R920 sensor_0.a.n0 sensor_0.a.t1 14.2976
R921 sensor_0.a sensor_0.a.n11 1.63801
R922 sensor_0.a.n11 sensor_0.a.n7 1.541
R923 sensor_0.a.n11 sensor_0.a.n10 1.541
R924 sensor_0.a.n10 sensor_0.a.n9 0.873387
R925 sensor_0.a.n6 sensor_0.a.n5 0.865287
R926 sensor_0.a.n7 sensor_0.a.n6 0.864262
R927 sensor_0.a.n9 sensor_0.a.n8 0.848309
R928 sensor_0.a.n3 sensor_0.a.n2 0.538
R929 sensor_0.a.n4 sensor_0.a.n3 0.538
R930 sensor_0.a.n0 sensor_0.a.n4 0.488
R931 sensor_0.a.n1 sensor_0.a.n0 0.29354
R932 sensor_0.a sensor_0.a.n1 0.28675
R933 vpwr.t13 vpwr.t26 790.188
R934 vpwr.t22 vpwr.t18 648.131
R935 vpwr.t4 vpwr.t10 583.023
R936 vpwr.n77 vpwr 548.548
R937 vpwr.n56 vpwr.t11 514.011
R938 vpwr.t8 vpwr.t22 485.358
R939 vpwr.t12 vpwr.t16 414.33
R940 vpwr.n14 vpwr.t3 413.315
R941 vpwr.n32 vpwr.t27 375.277
R942 vpwr.n7 vpwr.t0 344.005
R943 vpwr.t20 vpwr.t1 319.627
R944 vpwr.n50 vpwr.n39 311.957
R945 vpwr.n72 vpwr.n31 311.894
R946 vpwr.n59 vpwr.n58 309.18
R947 vpwr.t10 vpwr.t15 292.991
R948 vpwr.t24 vpwr.t12 292.991
R949 vpwr.n43 vpwr.n40 292.5
R950 vpwr.n45 vpwr.n44 292.5
R951 vpwr.t18 vpwr.t28 287.072
R952 vpwr.t16 vpwr.t4 287.072
R953 vpwr.t26 vpwr.t24 272.274
R954 vpwr.t15 vpwr.t25 254.518
R955 vpwr.t1 vpwr.t8 248.599
R956 vpwr.t25 vpwr.t20 248.599
R957 vpwr.t6 vpwr.t13 244.306
R958 vpwr.n6 vpwr.t31 187.321
R959 vpwr vpwr.t6 186.556
R960 vpwr.n44 vpwr.n43 182.929
R961 vpwr.n7 vpwr.n5 152
R962 vpwr.n42 vpwr.n41 148.689
R963 vpwr.n14 vpwr.t30 126.127
R964 vpwr.n39 vpwr.t21 119.608
R965 vpwr.n58 vpwr.t17 93.81
R966 vpwr.n6 vpwr.n1 73.2067
R967 vpwr.n43 vpwr.t9 68.0124
R968 vpwr.n58 vpwr.t5 63.3219
R969 vpwr.n39 vpwr.t2 63.3219
R970 vpwr.n41 vpwr.t19 61.9158
R971 vpwr.n31 vpwr.t14 41.5552
R972 vpwr.n31 vpwr.t7 41.5552
R973 vpwr.n71 vpwr.n70 34.6358
R974 vpwr.n64 vpwr.n34 34.6358
R975 vpwr.n65 vpwr.n64 34.6358
R976 vpwr.n66 vpwr.n65 34.6358
R977 vpwr.n60 vpwr.n57 34.6358
R978 vpwr.n51 vpwr.n37 34.6358
R979 vpwr.n55 vpwr.n37 34.6358
R980 vpwr.n66 vpwr.n32 32.377
R981 vpwr.n56 vpwr.n55 32.0005
R982 vpwr.n41 vpwr.t29 30.239
R983 vpwr.n50 vpwr.n49 30.1181
R984 vpwr.n44 vpwr.t23 29.316
R985 vpwr.n72 vpwr.n71 22.9652
R986 vpwr.n51 vpwr.n50 20.3299
R987 vpwr.n70 vpwr.n32 18.0711
R988 vpwr vpwr.n4 14.0185
R989 vpwr.n45 vpwr.n42 13.9946
R990 vpwr.n49 vpwr.n40 12.8758
R991 vpwr.n57 vpwr.n56 9.41227
R992 vpwr.n11 vpwr.n10 9.3005
R993 vpwr.n8 vpwr.n2 9.3005
R994 vpwr.n8 vpwr.n7 9.3005
R995 vpwr.n7 vpwr.n6 9.15991
R996 vpwr.n15 vpwr.n14 7.02651
R997 vpwr.n59 vpwr.n34 6.02403
R998 vpwr.n46 vpwr.n45 5.00414
R999 vpwr.n4 vpwr 4.7293
R1000 vpwr.n9 vpwr.n0 4.6505
R1001 vpwr.n18 vpwr.n17 4.6505
R1002 vpwr.n47 vpwr.n46 4.6505
R1003 vpwr.n49 vpwr.n48 4.6505
R1004 vpwr.n50 vpwr.n38 4.6505
R1005 vpwr.n52 vpwr.n51 4.6505
R1006 vpwr.n53 vpwr.n37 4.6505
R1007 vpwr.n55 vpwr.n54 4.6505
R1008 vpwr.n56 vpwr.n36 4.6505
R1009 vpwr.n57 vpwr.n35 4.6505
R1010 vpwr.n61 vpwr.n60 4.6505
R1011 vpwr.n62 vpwr.n34 4.6505
R1012 vpwr.n64 vpwr.n63 4.6505
R1013 vpwr.n65 vpwr.n33 4.6505
R1014 vpwr.n67 vpwr.n66 4.6505
R1015 vpwr.n68 vpwr.n32 4.6505
R1016 vpwr.n70 vpwr.n69 4.6505
R1017 vpwr.n71 vpwr.n30 4.6505
R1018 vpwr.n4 vpwr 4.53383
R1019 vpwr.n46 vpwr.n40 4.07323
R1020 vpwr.n73 vpwr.n72 3.93272
R1021 vpwr.n60 vpwr.n59 3.76521
R1022 vpwr.n5 vpwr 3.11401
R1023 vpwr.n17 vpwr.n15 3.0725
R1024 vpwr.n27 vpwr.n26 2.91783
R1025 vpwr.n28 vpwr 2.44425
R1026 vpwr.n12 vpwr 2.36657
R1027 vpwr.n5 vpwr.n1 1.55726
R1028 vpwr.n10 vpwr.n9 1.55726
R1029 vpwr.n8 vpwr.n1 1.38428
R1030 vpwr.n9 vpwr.n8 1.38428
R1031 vpwr.n10 vpwr 1.38428
R1032 vpwr.n17 vpwr.n16 1.2805
R1033 vpwr.n77 vpwr.n76 0.711611
R1034 vpwr.n12 vpwr 0.580857
R1035 vpwr.n29 vpwr.n28 0.5255
R1036 vpwr.n75 vpwr 0.223
R1037 vpwr.n3 vpwr 0.196446
R1038 vpwr.n20 vpwr 0.171696
R1039 vpwr.n47 vpwr.n42 0.144332
R1040 vpwr.n73 vpwr.n30 0.138831
R1041 vpwr.n48 vpwr.n47 0.120292
R1042 vpwr.n48 vpwr.n38 0.120292
R1043 vpwr.n52 vpwr.n38 0.120292
R1044 vpwr.n53 vpwr.n52 0.120292
R1045 vpwr.n54 vpwr.n53 0.120292
R1046 vpwr.n54 vpwr.n36 0.120292
R1047 vpwr.n36 vpwr.n35 0.120292
R1048 vpwr.n61 vpwr.n35 0.120292
R1049 vpwr.n62 vpwr.n61 0.120292
R1050 vpwr.n63 vpwr.n62 0.120292
R1051 vpwr.n63 vpwr.n33 0.120292
R1052 vpwr.n67 vpwr.n33 0.120292
R1053 vpwr.n68 vpwr.n67 0.120292
R1054 vpwr.n69 vpwr.n68 0.120292
R1055 vpwr.n69 vpwr.n30 0.120292
R1056 vpwr.n74 vpwr.n73 0.107496
R1057 vpwr.n20 vpwr.n19 0.0901739
R1058 vpwr vpwr.n83 0.0634013
R1059 vpwr.n27 vpwr 0.063
R1060 vpwr.n21 vpwr.n20 0.0500874
R1061 vpwr.n13 vpwr.n12 0.0466957
R1062 vpwr.n24 vpwr.n23 0.0435328
R1063 vpwr.n83 vpwr.n29 0.039096
R1064 vpwr.n18 vpwr.n13 0.0331087
R1065 vpwr.n83 vpwr.n82 0.0287348
R1066 vpwr.n3 vpwr.n2 0.02675
R1067 vpwr vpwr.n11 0.0255
R1068 vpwr.n22 vpwr.n21 0.0213989
R1069 vpwr.n78 vpwr.n75 0.0207266
R1070 vpwr.n26 vpwr.n25 0.018111
R1071 vpwr.n74 vpwr 0.0174271
R1072 vpwr vpwr.n74 0.01675
R1073 vpwr.n19 vpwr.n18 0.014087
R1074 vpwr.n24 vpwr.n22 0.0127951
R1075 vpwr.n11 vpwr.n0 0.01175
R1076 vpwr.n2 vpwr.n0 0.0105
R1077 vpwr.n81 vpwr.n80 0.009875
R1078 vpwr vpwr.n3 0.00725676
R1079 vpwr.n23 vpwr 0.00459836
R1080 vpwr.n79 vpwr.n78 0.00412592
R1081 vpwr.n80 vpwr.n79 0.003625
R1082 vpwr.n82 vpwr.n81 0.00196888
R1083 vpwr.n26 vpwr.n24 0.0016109
R1084 vpwr.n78 vpwr.n77 0.00154933
R1085 vpwr.n28 vpwr.n27 0.000500433
R1086 vtd.n7 vtd.t29 64.6821
R1087 vtd.n8 vtd.t27 64.3461
R1088 vtd.n4 vtd.t24 63.6317
R1089 vtd.n9 vtd.t26 63.6292
R1090 vtd.n8 vtd.t28 63.6292
R1091 vtd.n17 vtd.t18 63.6292
R1092 vtd.n2 vtd.t16 63.6292
R1093 vtd.n18 vtd.t14 63.6292
R1094 vtd.n1 vtd.t12 63.6292
R1095 vtd.n19 vtd.t20 63.6292
R1096 vtd.n0 vtd.t22 63.6292
R1097 vtd.n6 vtd.t8 63.6292
R1098 vtd.n3 vtd.t10 63.6275
R1099 vtd.n13 vtd.t4 18.2948
R1100 vtd.n10 vtd.t1 18.1899
R1101 vtd.n10 vtd.t5 17.4187
R1102 vtd.n13 vtd.t0 17.4177
R1103 vtd.n11 vtd.t2 17.4156
R1104 vtd.n14 vtd.t7 17.4136
R1105 vtd.n12 vtd.t6 17.4125
R1106 vtd.n15 vtd.t3 17.4115
R1107 vtd.n3 vtd.t11 14.3559
R1108 vtd.n17 vtd.t19 14.3555
R1109 vtd.n2 vtd.t15 14.283
R1110 vtd.n2 vtd.t17 14.283
R1111 vtd.n1 vtd.t21 14.283
R1112 vtd.n1 vtd.t13 14.283
R1113 vtd.n0 vtd.t9 14.283
R1114 vtd.n0 vtd.t23 14.283
R1115 vtd.n7 vtd.t25 13.7801
R1116 vtd.n16 vtd.n15 2.14635
R1117 vtd.n3 vtd.n16 1.54335
R1118 vtd vtd.n20 1.22372
R1119 vtd.n16 vtd.n12 1.09526
R1120 vtd.n20 vtd.n3 0.981002
R1121 vtd.n15 vtd.n14 0.8755
R1122 vtd.n14 vtd.n13 0.8755
R1123 vtd.n5 vtd.n7 0.832184
R1124 vtd.n11 vtd.n10 0.769433
R1125 vtd.n12 vtd.n11 0.769356
R1126 vtd.n9 vtd.n8 0.717388
R1127 vtd.n4 vtd.n9 0.708453
R1128 vtd.n20 vtd.n5 0.438348
R1129 vtd.n3 vtd.n6 0.140567
R1130 vtd.n18 vtd.n2 0.140142
R1131 vtd.n19 vtd.n1 0.140142
R1132 vtd.n6 vtd.n0 0.140142
R1133 vtd.n0 vtd.n19 0.134875
R1134 vtd.n1 vtd.n18 0.134875
R1135 vtd.n2 vtd.n17 0.134875
R1136 vtd.n5 vtd.n4 0.114328
R1137 vts.n33 vts.n27 7140
R1138 vts.n31 vts.n27 7140
R1139 vts.n31 vts.n26 6543.53
R1140 vts.n34 vts.n33 6017.65
R1141 vts.n29 vts.n28 761.601
R1142 vts.n30 vts.n29 761.601
R1143 vts.n30 vts.n25 697.977
R1144 vts.n28 vts.n23 641.883
R1145 vts.n37 vts.n26 596.471
R1146 vts.n34 vts.n24 592.942
R1147 vts.t7 vts.t22 338.649
R1148 vts.t4 vts.t18 333.303
R1149 vts.t22 vts.n27 262.014
R1150 vts.n35 vts.t18 237.054
R1151 vts.t2 vts.t4 229.925
R1152 vts.t0 vts.t2 229.925
R1153 vts.t15 vts.t0 229.925
R1154 vts.t13 vts.t11 229.925
R1155 vts.t11 vts.t9 229.925
R1156 vts.t9 vts.t7 229.925
R1157 vts.n32 vts.t15 130.113
R1158 vts.n32 vts.t13 99.8129
R1159 vts.n21 vts.t17 63.6292
R1160 vts.n14 vts.t21 63.6292
R1161 vts.n38 vts.n25 63.624
R1162 vts.n39 vts.n23 52.424
R1163 vts.n39 vts.n38 45.6476
R1164 vts.n1 vts.t31 27.6073
R1165 vts.n6 vts.t32 27.1628
R1166 vts.n5 vts.t25 26.7019
R1167 vts.n0 vts.t26 26.4053
R1168 vts.n0 vts.t34 26.2229
R1169 vts.n4 vts.t30 25.2012
R1170 vts.n2 vts.t33 25.2012
R1171 vts.n7 vts.t27 24.699
R1172 vts.n3 vts.t28 24.699
R1173 vts.n8 vts.t29 24.1526
R1174 vts.n42 vts.t6 16.8006
R1175 vts.n15 vts.t23 14.4639
R1176 vts.n20 vts.t20 14.4362
R1177 vts.n22 vts.t19 14.4313
R1178 vts.n14 vts.t24 14.3697
R1179 vts.n10 vts.t5 14.283
R1180 vts.n10 vts.t3 14.283
R1181 vts.n11 vts.t1 14.283
R1182 vts.n11 vts.t16 14.283
R1183 vts.n12 vts.t14 14.283
R1184 vts.n12 vts.t12 14.283
R1185 vts.n13 vts.t10 14.283
R1186 vts.n13 vts.t8 14.283
R1187 vts.n43 vts.n42 4.5005
R1188 vts.n44 vts 3.013
R1189 vts vts.n8 2.98635
R1190 vts.n5 vts.n4 2.30564
R1191 vts.n1 vts.n0 2.30482
R1192 vts.n3 vts.n2 2.27981
R1193 vts.n7 vts.n6 2.24388
R1194 vts vts.n44 2.01425
R1195 vts vts.n43 0.8255
R1196 vts.n6 vts.n5 0.680761
R1197 vts.n4 vts.n3 0.680308
R1198 vts.n8 vts.n7 0.680308
R1199 vts.n19 vts.n18 0.6455
R1200 vts.n18 vts.n17 0.6455
R1201 vts.n17 vts.n16 0.6455
R1202 vts.n2 vts.n1 0.604164
R1203 vts.n16 vts.n15 0.450361
R1204 vts.n20 vts.n19 0.440551
R1205 vts.n44 vts 0.26925
R1206 vts.n40 vts.n22 0.0947919
R1207 vts.n15 vts.n14 0.0741592
R1208 vts.n21 vts.n20 0.0682354
R1209 vts.n22 vts.n21 0.0634447
R1210 vts.n43 vts.n9 0.05093
R1211 vts.n34 vts.n23 0.0426316
R1212 vts.n35 vts.n34 0.0426316
R1213 vts.n26 vts.n25 0.0175052
R1214 vts.n35 vts.n26 0.0175052
R1215 vts.n19 vts.n10 0.0129196
R1216 vts.n18 vts.n11 0.0129196
R1217 vts.n17 vts.n12 0.0129196
R1218 vts.n16 vts.n13 0.0129196
R1219 vts.n37 vts.n36 0.011183
R1220 vts.n38 vts.n37 0.0106833
R1221 vts.n36 vts.n24 0.0075124
R1222 vts.n39 vts.n9 0.00749235
R1223 vts.n39 vts.n24 0.00701261
R1224 vts.n29 vts.n27 0.00559165
R1225 vts.n33 vts.n28 0.00192573
R1226 vts.n33 vts.n32 0.00192573
R1227 vts.n31 vts.n30 0.00192573
R1228 vts.n32 vts.n31 0.00192573
R1229 vts.n41 vts.n9 0.00151802
R1230 vts.n41 vts.n40 0.00150795
R1231 vts.n36 vts.n35 0.00100013
R1232 vts.n40 vts.n39 0.00100001
R1233 vts.n42 vts.n41 0.001
R1234 buffer_0.b.n0 buffer_0.b.t11 40.2461
R1235 buffer_0.b.n2 buffer_0.b.t10 40.2461
R1236 buffer_0.b buffer_0.b.t9 39.5317
R1237 buffer_0.b.n1 buffer_0.b.t16 39.5292
R1238 buffer_0.b.n1 buffer_0.b.t18 39.5292
R1239 buffer_0.b.n0 buffer_0.b.t13 39.5292
R1240 buffer_0.b.n0 buffer_0.b.t14 39.5292
R1241 buffer_0.b.n3 buffer_0.b.t12 39.5292
R1242 buffer_0.b.n3 buffer_0.b.t19 39.5292
R1243 buffer_0.b.n2 buffer_0.b.t17 39.5292
R1244 buffer_0.b.n2 buffer_0.b.t15 39.5292
R1245 buffer_0.b.n4 buffer_0.b.t6 17.4005
R1246 buffer_0.b.n4 buffer_0.b.t2 17.4005
R1247 buffer_0.b.n5 buffer_0.b.t4 17.4005
R1248 buffer_0.b.n5 buffer_0.b.t7 17.4005
R1249 buffer_0.b.n6 buffer_0.b.t3 17.4005
R1250 buffer_0.b.n6 buffer_0.b.t8 17.4005
R1251 buffer_0.b.n7 buffer_0.b.t5 17.4005
R1252 buffer_0.b.n7 buffer_0.b.t1 17.4005
R1253 buffer_0.b.n4 buffer_0.b.n5 3.17349
R1254 buffer_0.b.n6 buffer_0.b.n7 2.69321
R1255 buffer_0.b.n5 buffer_0.b.n6 2.68836
R1256 buffer_0.b.t0 buffer_0.b.n4 2.65092
R1257 buffer_0.b.n3 buffer_0.b.n2 2.15117
R1258 buffer_0.b.n1 buffer_0.b.n0 2.15117
R1259 buffer_0.b buffer_0.b.n1 1.49152
R1260 buffer_0.b buffer_0.b.t0 0.968485
R1261 buffer_0.b buffer_0.b.n3 0.961845
R1262 buffer_0.c buffer_0.c.t10 18.4486
R1263 buffer_0.c.n17 buffer_0.c.t16 17.4005
R1264 buffer_0.c.n17 buffer_0.c.t6 17.4005
R1265 buffer_0.c.n15 buffer_0.c.t7 17.4005
R1266 buffer_0.c.n15 buffer_0.c.t18 17.4005
R1267 buffer_0.c.n13 buffer_0.c.t13 17.4005
R1268 buffer_0.c.n13 buffer_0.c.t1 17.4005
R1269 buffer_0.c.n11 buffer_0.c.t2 17.4005
R1270 buffer_0.c.n11 buffer_0.c.t20 17.4005
R1271 buffer_0.c.n7 buffer_0.c.t4 17.4005
R1272 buffer_0.c.n7 buffer_0.c.t17 17.4005
R1273 buffer_0.c.n5 buffer_0.c.t12 17.4005
R1274 buffer_0.c.n5 buffer_0.c.t3 17.4005
R1275 buffer_0.c.n3 buffer_0.c.t0 17.4005
R1276 buffer_0.c.n3 buffer_0.c.t14 17.4005
R1277 buffer_0.c.n1 buffer_0.c.t11 17.4005
R1278 buffer_0.c.n1 buffer_0.c.t8 17.4005
R1279 buffer_0.c.n0 buffer_0.c.t5 17.4005
R1280 buffer_0.c.n0 buffer_0.c.t19 17.4005
R1281 buffer_0.c.n9 buffer_0.c.t15 17.4005
R1282 buffer_0.c.n9 buffer_0.c.t9 17.4005
R1283 buffer_0.c.n2 buffer_0.c.n0 1.87829
R1284 buffer_0.c buffer_0.c.n18 1.52139
R1285 buffer_0.c.n18 buffer_0.c.n17 1.51465
R1286 buffer_0.c.n4 buffer_0.c.n2 1.08383
R1287 buffer_0.c.n6 buffer_0.c.n4 1.08383
R1288 buffer_0.c.n10 buffer_0.c.n8 1.08383
R1289 buffer_0.c.n12 buffer_0.c.n10 1.08383
R1290 buffer_0.c.n14 buffer_0.c.n12 1.08383
R1291 buffer_0.c.n8 buffer_0.c.n6 1.04217
R1292 buffer_0.c.n16 buffer_0.c.n14 1.04217
R1293 buffer_0.c.n6 buffer_0.c.n5 0.776026
R1294 buffer_0.c.n14 buffer_0.c.n13 0.766495
R1295 buffer_0.c.n4 buffer_0.c.n3 0.766495
R1296 buffer_0.c.n16 buffer_0.c.n15 0.766495
R1297 buffer_0.c.n12 buffer_0.c.n11 0.766495
R1298 buffer_0.c.n8 buffer_0.c.n7 0.766495
R1299 buffer_0.c.n2 buffer_0.c.n1 0.766495
R1300 buffer_0.c.n10 buffer_0.c.n9 0.766495
R1301 buffer_0.c.n18 buffer_0.c.n16 0.333833
R1302 ib.n1 ib.t5 38.0465
R1303 ib.n1 ib.t0 37.3602
R1304 ib.n3 ib.t2 18.7313
R1305 ib.n3 ib.t4 17.409
R1306 ib.n0 ib.t1 17.4005
R1307 ib.n0 ib.t3 17.4005
R1308 ib ib.n4 1.76488
R1309 ib.n2 ib.n1 0.239515
R1310 ib.n4 ib.n3 0.0163842
R1311 ib.n2 ib.n0 0.00444823
R1312 ib.n4 ib.n2 0.00358796
R1313 out_sigma.n1 out_sigma.t2 394.808
R1314 out_sigma.n0 out_sigma.t0 250.941
R1315 out_sigma out_sigma.t1 144.601
R1316 out_sigma out_sigma.n1 9.0826
R1317 out_sigma out_sigma.n0 4.7225
R1318 out_sigma.n2 out_sigma 3.8755
R1319 out_sigma.n0 out_sigma 3.35288
R1320 out_sigma.n2 out_sigma 3.2272
R1321 out_sigma.n1 out_sigma 0.727062
R1322 out_sigma out_sigma.n2 0.13175
R1323 clk.n0 clk.t0 294.557
R1324 clk.n0 clk.t1 211.01
R1325 clk.n2 clk.n0 8.28655
R1326 clk.n3 clk 7.73487
R1327 clk.n3 clk.n2 1.82961
R1328 clk.n1 clk 0.981259
R1329 clk.n2 clk.n1 0.848973
R1330 clk clk.n5 0.385917
R1331 clk.n5 clk.n4 0.03175
R1332 clk.n4 clk.n3 0.00111796
R1333 out.n2 out.t0 8.97158
R1334 out.n2 out.n1 2.56714
R1335 out.n0 out.t2 0.506271
R1336 out.n1 out.n0 0.504061
R1337 out out.n2 0.240344
R1338 out.n0 out.t1 0.0277714
R1339 out.n1 out.t3 0.00303875
C0 buffer_0.d buffer_0.b 1.04f
C1 buffer_0.a ib 0.0615f
C2 a_15712_3988# a_16854_3988# 0.00957f
C3 a_15048_3988# vd 0.00206f
C4 vts ib 2.21f
C5 a_16854_3988# sigma-delta_0.x1.D 2.69e-19
C6 a_16190_3988# out_buff 9.87e-22
C7 a_16190_3988# a_15712_3988# 0.357f
C8 a_16522_3988# vpwr 0.00266f
C9 out out_buff 0.0112f
C10 a_15712_3988# out 0.18f
C11 vd vpwr 0.00726f
C12 a_17020_5320# sigma-delta_0.x1.Q 0.00839f
C13 a_14550_5320# out_sigma 6.23e-19
C14 buffer_0.c out 8.56e-19
C15 a_15881_2489# a_15706_2515# 0.251f
C16 sensor_0.c sensor_0.b 0.55f
C17 a_15359_2757# a_15141_2515# 0.21f
C18 a_16356_5320# a_16024_5320# 0.3f
C19 buffer_0.b ib 0.0167f
C20 vd a_16522_3988# 0.00558f
C21 a_15881_2489# clk 2.68e-20
C22 a_15881_2489# a_15712_3988# 0.00381f
C23 a_15706_2515# a_15141_2515# 7.99e-20
C24 a_15881_2489# sigma-delta_0.x1.D 0.004f
C25 a_15359_2757# sigma-delta_0.x1.Q 0.00111f
C26 vpwr a_16060_2515# 0.00312f
C27 clk a_15141_2515# 3.26e-19
C28 vts sensor_0.b 1f
C29 a_15712_3988# a_15141_2515# 2.02e-20
C30 a_15881_2489# a_14625_2515# 0.0436f
C31 a_15706_2515# sigma-delta_0.x1.Q 0.00593f
C32 a_15141_2515# sigma-delta_0.x1.D 0.00353f
C33 a_15359_2757# a_14791_2515# 0.186f
C34 a_16190_3988# vpwr 0.00384f
C35 a_15380_3988# a_15141_2515# 1.22e-19
C36 a_14716_3988# a_14882_5320# 0.00434f
C37 buffer_0.d ib 0.194f
C38 a_15712_3988# sigma-delta_0.x1.Q 0.414f
C39 a_15706_2515# a_14791_2515# 0.125f
C40 a_14882_5320# out_buff 0.0014f
C41 a_15141_2515# a_14625_2515# 0.115f
C42 sigma-delta_0.x1.D sigma-delta_0.x1.Q 0.0675f
C43 out_sigma a_15359_2757# 3.73e-19
C44 buffer_0.a out_buff 3.96f
C45 a_16854_3988# a_16522_3988# 0.303f
C46 a_16024_5320# out_buff 3.49e-20
C47 a_15712_3988# a_16024_5320# 0.00827f
C48 a_15380_3988# sigma-delta_0.x1.Q 1.43e-21
C49 vts out_buff 2.36f
C50 clk a_14791_2515# 0.00241f
C51 a_14791_2515# out_buff 8.29e-20
C52 a_15712_3988# a_14791_2515# 4.13e-19
C53 a_16190_3988# a_16522_3988# 0.312f
C54 a_15706_2515# out_sigma 6.85e-19
C55 buffer_0.a buffer_0.c 3.88f
C56 vd a_16854_3988# 0.0174f
C57 sigma-delta_0.x1.Q a_14625_2515# 9.54e-19
C58 a_15712_3988# a_15546_5320# 0.00466f
C59 a_15546_5320# out_buff 2.84e-19
C60 sigma-delta_0.x1.D a_14791_2515# 0.229f
C61 vts buffer_0.c 1.08f
C62 out_sigma a_14716_3988# 0.0146f
C63 a_15359_2757# a_15237_2515# 3.16e-19
C64 a_16190_3988# vd 0.00388f
C65 a_15706_2515# a_16445_2515# 7.05e-19
C66 a_15881_2489# vpwr 0.688f
C67 out_sigma clk 0.382f
C68 vd out 0.145p
C69 out_sigma out_buff 2.19f
C70 a_15380_3988# a_15546_5320# 0.00434f
C71 a_15868_2881# a_15359_2757# 2.6e-19
C72 a_15712_3988# out_sigma 0.16f
C73 a_15249_2881# a_15141_2515# 0.0572f
C74 a_14791_2515# a_14625_2515# 0.906f
C75 out_sigma sigma-delta_0.x1.D 0.294f
C76 a_17020_5320# a_16688_5320# 0.299f
C77 a_15712_3988# a_16445_2515# 0.00366f
C78 a_15380_3988# out_sigma 0.0148f
C79 out_sigma buffer_0.c 0.00107f
C80 vd sensor_0.a 2.92f
C81 a_15868_2881# a_15706_2515# 0.00645f
C82 a_15046_2515# a_15141_2515# 0.0498f
C83 a_16445_2515# sigma-delta_0.x1.D 0.00209f
C84 a_16356_5320# a_16688_5320# 0.307f
C85 a_15249_2881# sigma-delta_0.x1.Q 3.66e-19
C86 buffer_0.b out_buff 2.8f
C87 a_15141_2515# vpwr 0.363f
C88 clk a_15237_2515# 5.33e-20
C89 out_sigma a_14625_2515# 0.00261f
C90 a_15048_3988# a_14882_5320# 0.00482f
C91 a_15881_2489# a_16522_3988# 1.28e-20
C92 a_15141_2515# a_15403_2515# 0.00171f
C93 a_15868_2881# a_15712_3988# 5.54e-20
C94 sigma-delta_0.x1.D a_15237_2515# 8.22e-19
C95 buffer_0.b buffer_0.c 1.34f
C96 a_15214_5320# out_buff 5.44e-19
C97 a_16445_2515# a_14625_2515# 4.71e-20
C98 a_15046_2515# sigma-delta_0.x1.Q 7.58e-20
C99 a_15881_2489# vd 0.00172f
C100 a_15868_2881# sigma-delta_0.x1.D 2.11e-20
C101 a_15249_2881# a_14791_2515# 0.0346f
C102 vpwr sigma-delta_0.x1.Q 0.186f
C103 a_15048_3988# a_14791_2515# 1.82e-19
C104 sensor_0.b sensor_0.d 0.0152f
C105 a_15214_5320# a_15380_3988# 0.00473f
C106 sigma-delta_0.x1.Q a_15403_2515# 9.75e-20
C107 a_14625_2515# a_15237_2515# 0.00134f
C108 a_15046_2515# a_14791_2515# 0.0642f
C109 a_14791_2515# vpwr 0.607f
C110 a_15048_3988# out_sigma 0.0146f
C111 vd sensor_0.c 0.804f
C112 buffer_0.d clk 0.202f
C113 buffer_0.d out_buff 40.1f
C114 vd a_6126_29386# 0.0189f
C115 a_15359_2757# a_15815_2515# 4.2e-19
C116 a_16522_3988# sigma-delta_0.x1.Q 5e-20
C117 buffer_0.d buffer_0.c 1.32f
C118 ib sensor_0.b 2.02e-19
C119 out_sigma vpwr 2.04f
C120 vd sigma-delta_0.x1.Q 0.0969f
C121 a_15712_3988# a_16688_5320# 0.00557f
C122 a_15706_2515# a_15815_2515# 0.00742f
C123 a_15881_2489# a_16060_2515# 0.0074f
C124 vd a_14882_5320# 0.061f
C125 vd buffer_0.a 6.66f
C126 a_16445_2515# vpwr 0.2f
C127 a_16024_5320# vd 0.0626f
C128 a_15048_3988# a_15214_5320# 0.00473f
C129 vts vd 1.62f
C130 clk a_15815_2515# 1.1e-20
C131 a_15046_2515# a_15237_2515# 4.61e-19
C132 vd a_14791_2515# 1.08e-19
C133 a_15712_3988# a_15815_2515# 1.36e-20
C134 a_15881_2489# a_16190_3988# 4.27e-19
C135 vpwr a_15237_2515# 0.00292f
C136 a_14550_5320# a_14716_3988# 0.00458f
C137 a_15546_5320# vd 0.0619f
C138 sigma-delta_0.x1.D a_15815_2515# 2.42e-20
C139 a_15868_2881# vpwr 9.63e-19
C140 a_14550_5320# out_buff 0.0535f
C141 ib out_buff 0.0112f
C142 vd out_sigma 1.88f
C143 a_16445_2515# a_16522_3988# 1.4e-19
C144 a_16060_2515# sigma-delta_0.x1.Q 6.05e-19
C145 a_15815_2515# a_14625_2515# 2.56e-19
C146 ib buffer_0.c 0.0951f
C147 vd a_16445_2515# 0.00317f
C148 a_6126_29386# out 0.0171f
C149 a_16854_3988# sigma-delta_0.x1.Q 0.414f
C150 vd buffer_0.b 6.37f
C151 a_16190_3988# sigma-delta_0.x1.Q 1.87e-20
C152 sensor_0.a sensor_0.c 0.997f
C153 a_15712_3988# a_17020_5320# 0.00974f
C154 a_15214_5320# vd 0.0598f
C155 a_14882_5320# out 0.0019f
C156 a_16356_5320# a_15712_3988# 0.00631f
C157 a_16190_3988# a_16024_5320# 0.00473f
C158 buffer_0.a out 0.0533f
C159 a_16024_5320# out 0.00189f
C160 vts out 0.00336f
C161 a_15706_2515# a_15359_2757# 0.0512f
C162 a_16854_3988# out_sigma 7.61e-19
C163 a_15546_5320# out 0.00187f
C164 vpwr a_15815_2515# 7.93e-19
C165 vts sensor_0.a 0.543f
C166 buffer_0.d vd 2.79f
C167 clk a_15359_2757# 1.78e-19
C168 a_15712_3988# a_15359_2757# 7.49e-21
C169 a_16522_3988# a_16688_5320# 0.00482f
C170 a_15881_2489# sigma-delta_0.x1.Q 0.142f
C171 out_sigma out 5.44f
C172 a_15359_2757# sigma-delta_0.x1.D 6.24e-19
C173 vd a_16688_5320# 0.0633f
C174 a_15706_2515# clk 6.46e-20
C175 vd sensor_0.d 0.282f
C176 a_15380_3988# a_15359_2757# 7.2e-20
C177 a_15706_2515# a_15712_3988# 0.0011f
C178 buffer_0.b out 0.0634f
C179 a_15881_2489# a_14791_2515# 0.0426f
C180 a_15706_2515# sigma-delta_0.x1.D 9.45e-19
C181 a_15712_3988# a_14716_3988# 2.04e-19
C182 a_14716_3988# out_buff 0.307f
C183 a_15141_2515# sigma-delta_0.x1.Q 8.11e-19
C184 a_15359_2757# a_14625_2515# 0.0701f
C185 clk out_buff 0.843f
C186 sigma-delta_0.x1.D a_14716_3988# 2.07e-19
C187 a_15712_3988# out_buff 0.00915f
C188 a_15214_5320# out 0.00184f
C189 clk sigma-delta_0.x1.D 0.00993f
C190 sigma-delta_0.x1.D out_buff 1.65e-19
C191 a_15712_3988# sigma-delta_0.x1.D 0.339f
C192 a_15706_2515# a_14625_2515# 0.102f
C193 a_15881_2489# out_sigma 0.00735f
C194 vts sensor_0.c 0.192f
C195 a_14550_5320# vd 0.067f
C196 vd ib 0.0605f
C197 a_15141_2515# a_14791_2515# 0.23f
C198 buffer_0.c out_buff 2.02f
C199 a_15712_3988# a_15380_3988# 0.298f
C200 a_15380_3988# out_buff 5.35e-19
C201 a_14716_3988# a_14625_2515# 1.47e-19
C202 a_15881_2489# a_16445_2515# 0.107f
C203 clk a_14625_2515# 0.274f
C204 a_14625_2515# out_buff 4.76e-19
C205 a_15712_3988# a_14625_2515# 1.78e-19
C206 a_15249_2881# a_15359_2757# 0.0977f
C207 sigma-delta_0.x1.D a_14625_2515# 0.195f
C208 a_14791_2515# sigma-delta_0.x1.Q 0.00137f
C209 out_sigma a_15141_2515# 7.05e-19
C210 buffer_0.d out 0.00472f
C211 a_16854_3988# a_16688_5320# 0.00473f
C212 vts buffer_0.a 0.658f
C213 a_16356_5320# a_16522_3988# 0.00509f
C214 a_15359_2757# vpwr 0.378f
C215 vd a_17020_5320# 0.201f
C216 a_16024_5320# a_15546_5320# 0.144f
C217 out_sigma sigma-delta_0.x1.Q 0.668f
C218 a_16688_5320# out 0.00185f
C219 a_15048_3988# a_14716_3988# 0.296f
C220 a_16356_5320# vd 0.0637f
C221 a_15359_2757# a_15403_2515# 3.69e-19
C222 a_15141_2515# a_15237_2515# 0.0138f
C223 a_15048_3988# a_15712_3988# 4.38e-19
C224 a_15048_3988# out_buff 0.00138f
C225 buffer_0.a out_sigma 0.0172f
C226 a_15706_2515# vpwr 0.524f
C227 a_16445_2515# sigma-delta_0.x1.Q 0.226f
C228 a_15249_2881# sigma-delta_0.x1.D 5.56e-20
C229 sensor_0.a sensor_0.d 0.588f
C230 a_15048_3988# sigma-delta_0.x1.D 2.56e-20
C231 vts out_sigma 0.0608f
C232 out_sigma a_14791_2515# 0.00128f
C233 a_14716_3988# vpwr 0.0038f
C234 clk a_15046_2515# 3.09e-19
C235 a_15048_3988# a_15380_3988# 0.302f
C236 sigma-delta_0.x1.Q a_15237_2515# 1.45e-19
C237 clk vpwr 0.493f
C238 a_15712_3988# vpwr 0.0132f
C239 vpwr out_buff 0.0121f
C240 buffer_0.a buffer_0.b 0.126f
C241 a_15046_2515# sigma-delta_0.x1.D 0.164f
C242 a_16445_2515# a_14791_2515# 2.01e-19
C243 a_14550_5320# out 0.00197f
C244 a_15249_2881# a_14625_2515# 9.73e-19
C245 a_15868_2881# sigma-delta_0.x1.Q 4.53e-20
C246 vd sensor_0.b 0.0693f
C247 a_15048_3988# a_14625_2515# 1.92e-19
C248 sigma-delta_0.x1.D vpwr 0.483f
C249 clk a_15403_2515# 1.82e-20
C250 vts buffer_0.b 2.94f
C251 a_15214_5320# a_14882_5320# 0.303f
C252 a_15380_3988# vpwr 0.00397f
C253 a_14791_2515# a_15237_2515# 2.28e-19
C254 sigma-delta_0.x1.D a_15403_2515# 5.41e-20
C255 a_15046_2515# a_14625_2515# 0.0931f
C256 out_sigma a_16445_2515# 0.0691f
C257 a_15706_2515# vd 3.52e-19
C258 a_15868_2881# a_14791_2515# 1.46e-19
C259 vpwr a_14625_2515# 0.772f
C260 a_16854_3988# a_17020_5320# 0.00434f
C261 a_15712_3988# a_16522_3988# 0.0502f
C262 buffer_0.b out_sigma 0.017f
C263 vd a_14716_3988# 0.0021f
C264 a_15214_5320# a_15546_5320# 0.296f
C265 sensor_0.c sensor_0.d 0.492f
C266 a_17020_5320# out 0.00192f
C267 vd out_buff 3.22f
C268 a_15712_3988# vd 0.75f
C269 a_16190_3988# a_16356_5320# 0.00536f
C270 buffer_0.d buffer_0.a 2.4f
C271 vd sigma-delta_0.x1.D 0.908f
C272 a_16356_5320# out 0.00195f
C273 vts buffer_0.d 0.255f
C274 a_15380_3988# vd 0.00209f
C275 vd buffer_0.c 0.399f
C276 a_16688_5320# sigma-delta_0.x1.Q 0.0032f
C277 a_15249_2881# vpwr 0.156f
C278 a_15048_3988# vpwr 0.00379f
C279 vd a_14625_2515# 1.72e-20
C280 sensor_0.c ib 0.00238f
C281 vts sensor_0.d 0.248f
C282 a_15815_2515# sigma-delta_0.x1.Q 1.47e-19
C283 buffer_0.d out_sigma 0.0558f
C284 a_15046_2515# vpwr 0.0861f
C285 clk a_16060_2515# 6.32e-21
C286 vpwr a_15403_2515# 0.00407f
C287 a_14550_5320# a_14882_5320# 0.296f
C288 sensor_0.a sensor_0.b 0.821f
C289 a_14791_2515# a_15815_2515# 2.36e-20
C290 sigma-delta_0.x1.D a_16060_2515# 4.54e-20
C291 clk gnd 3.22f
C292 ib gnd 7.61f
C293 out_buff gnd 17.6f
C294 out gnd 59.7f
C295 out_sigma gnd 18.2f
C296 vpwr gnd 7.04f
C297 vts gnd 24.6f
C298 vd gnd 77.8f
C299 a_16060_2515# gnd 0.00223f
C300 a_15815_2515# gnd 9.68e-19
C301 a_15403_2515# gnd 0.00579f
C302 a_15237_2515# gnd 0.00863f
C303 a_15249_2881# gnd 0.00469f
C304 a_15046_2515# gnd 0.08f
C305 a_16445_2515# gnd 0.213f
C306 a_15706_2515# gnd 0.275f
C307 a_15881_2489# gnd 0.74f
C308 a_15141_2515# gnd 0.281f
C309 a_15359_2757# gnd 0.194f
C310 a_14791_2515# gnd 0.332f
C311 sigma-delta_0.x1.D gnd 2.56f
C312 a_14625_2515# gnd 0.7f
C313 sigma-delta_0.x1.Q gnd 1.09f
C314 a_17020_5320# gnd 0.557f
C315 a_16854_3988# gnd 0.348f
C316 a_16688_5320# gnd 0.388f
C317 a_16522_3988# gnd 0.356f
C318 a_16356_5320# gnd 0.392f
C319 a_16190_3988# gnd 0.357f
C320 a_16024_5320# gnd 0.447f
C321 a_15712_3988# gnd 69.7f
C322 a_15546_5320# gnd 0.449f
C323 a_15380_3988# gnd 0.365f
C324 a_15214_5320# gnd 0.387f
C325 a_15048_3988# gnd 0.364f
C326 a_14882_5320# gnd 0.39f
C327 a_14716_3988# gnd 0.366f
C328 buffer_0.c gnd 2.18f
C329 sensor_0.b gnd 16.7f
C330 sensor_0.c gnd 0.658f
C331 sensor_0.a gnd 5.59f
C332 sensor_0.d gnd 0.293f
C333 a_14550_5320# gnd 0.587f
C334 buffer_0.d gnd 27.6f
C335 buffer_0.b gnd 4.08f
C336 buffer_0.a gnd 5.13f
C337 a_6126_29386# gnd 0.593f
C338 out.t0 gnd 0.00791f
C339 out.t3 gnd 13.1f
C340 out.t2 gnd 29f
C341 out.t1 gnd 19.9f
C342 out.n0 gnd 10.6f
C343 out.n1 gnd 16.3f
C344 out.n2 gnd 61.5f
C345 out_sigma.t0 gnd 0.0145f
C346 out_sigma.t1 gnd 0.0107f
C347 out_sigma.n0 gnd 0.237f
C348 out_sigma.t2 gnd 0.0315f
C349 out_sigma.n1 gnd 2.76f
C350 out_sigma.n2 gnd 1.61f
C351 ib.t1 gnd 0.00293f
C352 ib.t3 gnd 0.00293f
C353 ib.n0 gnd 0.00778f
C354 ib.t5 gnd 0.0701f
C355 ib.t0 gnd 0.0693f
C356 ib.n1 gnd 0.0831f
C357 ib.n2 gnd 0.0236f
C358 ib.t4 gnd 0.00295f
C359 ib.t2 gnd 0.0315f
C360 ib.n3 gnd 0.139f
C361 ib.n4 gnd 0.0491f
C362 buffer_0.c.t5 gnd 0.0162f
C363 buffer_0.c.t19 gnd 0.0162f
C364 buffer_0.c.n0 gnd 0.356f
C365 buffer_0.c.t11 gnd 0.0162f
C366 buffer_0.c.t8 gnd 0.0162f
C367 buffer_0.c.n1 gnd 0.258f
C368 buffer_0.c.n2 gnd 0.326f
C369 buffer_0.c.t0 gnd 0.0162f
C370 buffer_0.c.t14 gnd 0.0162f
C371 buffer_0.c.n3 gnd 0.258f
C372 buffer_0.c.n4 gnd 0.25f
C373 buffer_0.c.t12 gnd 0.0162f
C374 buffer_0.c.t3 gnd 0.0162f
C375 buffer_0.c.n5 gnd 0.257f
C376 buffer_0.c.n6 gnd 0.249f
C377 buffer_0.c.t4 gnd 0.0162f
C378 buffer_0.c.t17 gnd 0.0162f
C379 buffer_0.c.n7 gnd 0.258f
C380 buffer_0.c.n8 gnd 0.247f
C381 buffer_0.c.t15 gnd 0.0162f
C382 buffer_0.c.t9 gnd 0.0162f
C383 buffer_0.c.n9 gnd 0.259f
C384 buffer_0.c.n10 gnd 0.25f
C385 buffer_0.c.t2 gnd 0.0162f
C386 buffer_0.c.t20 gnd 0.0162f
C387 buffer_0.c.n11 gnd 0.258f
C388 buffer_0.c.n12 gnd 0.25f
C389 buffer_0.c.t13 gnd 0.0162f
C390 buffer_0.c.t1 gnd 0.0162f
C391 buffer_0.c.n13 gnd 0.258f
C392 buffer_0.c.n14 gnd 0.247f
C393 buffer_0.c.t7 gnd 0.0162f
C394 buffer_0.c.t18 gnd 0.0162f
C395 buffer_0.c.n15 gnd 0.258f
C396 buffer_0.c.n16 gnd 0.187f
C397 buffer_0.c.t16 gnd 0.0162f
C398 buffer_0.c.t6 gnd 0.0162f
C399 buffer_0.c.n17 gnd 0.333f
C400 buffer_0.c.n18 gnd 0.298f
C401 buffer_0.c.t10 gnd 0.0328f
C402 buffer_0.b.n0 gnd 0.787f
C403 buffer_0.b.n1 gnd 0.539f
C404 buffer_0.b.n2 gnd 0.787f
C405 buffer_0.b.n3 gnd 0.619f
C406 buffer_0.b.n4 gnd 0.789f
C407 buffer_0.b.n5 gnd 0.719f
C408 buffer_0.b.n6 gnd 0.798f
C409 buffer_0.b.t10 gnd 0.465f
C410 buffer_0.b.t15 gnd 0.46f
C411 buffer_0.b.t17 gnd 0.46f
C412 buffer_0.b.t19 gnd 0.46f
C413 buffer_0.b.t12 gnd 0.46f
C414 buffer_0.b.t9 gnd 0.46f
C415 buffer_0.b.t16 gnd 0.46f
C416 buffer_0.b.t18 gnd 0.46f
C417 buffer_0.b.t13 gnd 0.46f
C418 buffer_0.b.t14 gnd 0.46f
C419 buffer_0.b.t11 gnd 0.465f
C420 buffer_0.b.t6 gnd 0.0187f
C421 buffer_0.b.t2 gnd 0.0187f
C422 buffer_0.b.t4 gnd 0.0187f
C423 buffer_0.b.t7 gnd 0.0187f
C424 buffer_0.b.t3 gnd 0.0187f
C425 buffer_0.b.t8 gnd 0.0187f
C426 buffer_0.b.t5 gnd 0.0187f
C427 buffer_0.b.t1 gnd 0.0187f
C428 buffer_0.b.n7 gnd 0.505f
C429 buffer_0.b.t0 gnd 0.607f
C430 vts.t26 gnd 0.102f
C431 vts.t34 gnd 0.101f
C432 vts.n0 gnd 0.158f
C433 vts.t31 gnd 0.103f
C434 vts.n1 gnd 0.0959f
C435 vts.t33 gnd 0.099f
C436 vts.n2 gnd 0.103f
C437 vts.t28 gnd 0.098f
C438 vts.n3 gnd 0.103f
C439 vts.t30 gnd 0.099f
C440 vts.n4 gnd 0.101f
C441 vts.t25 gnd 0.102f
C442 vts.n5 gnd 0.0979f
C443 vts.t32 gnd 0.103f
C444 vts.n6 gnd 0.0975f
C445 vts.t27 gnd 0.098f
C446 vts.n7 gnd 0.103f
C447 vts.t29 gnd 0.0968f
C448 vts.n8 gnd 0.147f
C449 vts.n9 gnd 0.0036f
C450 vts.t6 gnd 0.0681f
C451 vts.t17 gnd 0.18f
C452 vts.t20 gnd 0.011f
C453 vts.t5 gnd 0.0103f
C454 vts.t3 gnd 0.0103f
C455 vts.n10 gnd 0.0489f
C456 vts.t1 gnd 0.0103f
C457 vts.t16 gnd 0.0103f
C458 vts.n11 gnd 0.0489f
C459 vts.t14 gnd 0.0103f
C460 vts.t12 gnd 0.0103f
C461 vts.n12 gnd 0.0489f
C462 vts.t10 gnd 0.0103f
C463 vts.t8 gnd 0.0103f
C464 vts.n13 gnd 0.0489f
C465 vts.t23 gnd 0.0111f
C466 vts.t21 gnd 0.18f
C467 vts.t24 gnd 0.0108f
C468 vts.n14 gnd 0.216f
C469 vts.n15 gnd 0.123f
C470 vts.n16 gnd 0.0829f
C471 vts.n17 gnd 0.0968f
C472 vts.n18 gnd 0.0968f
C473 vts.n19 gnd 0.0822f
C474 vts.n20 gnd 0.123f
C475 vts.n21 gnd 0.116f
C476 vts.t19 gnd 0.011f
C477 vts.n22 gnd 0.0986f
C478 vts.n23 gnd 0.0571f
C479 vts.n24 gnd 0.00961f
C480 vts.n25 gnd 0.062f
C481 vts.n26 gnd 0.062f
C482 vts.t18 gnd 0.606f
C483 vts.n27 gnd 0.503f
C484 vts.n28 gnd 0.113f
C485 vts.t4 gnd 0.599f
C486 vts.t2 gnd 0.489f
C487 vts.t0 gnd 0.489f
C488 vts.t15 gnd 0.383f
C489 vts.t22 gnd 0.638f
C490 vts.t7 gnd 0.604f
C491 vts.t9 gnd 0.489f
C492 vts.t11 gnd 0.489f
C493 vts.t13 gnd 0.35f
C494 vts.n29 gnd 0.124f
C495 vts.n30 gnd 0.118f
C496 vts.n31 gnd 0.118f
C497 vts.n32 gnd 0.244f
C498 vts.n33 gnd 0.113f
C499 vts.n34 gnd 0.0575f
C500 vts.n35 gnd 0.352f
C501 vts.n37 gnd 0.00964f
C502 vts.n38 gnd 0.00928f
C503 vts.n39 gnd 0.0186f
C504 vts.n40 gnd 0.00808f
C505 vts.n41 gnd 0.00148f
C506 vts.n42 gnd 0.615f
C507 vts.n43 gnd 0.0622f
C508 vts.n44 gnd 1.57f
C509 vtd.n0 gnd 0.548f
C510 vtd.n1 gnd 0.548f
C511 vtd.n2 gnd 0.548f
C512 vtd.n3 gnd 0.963f
C513 vtd.n4 gnd 0.175f
C514 vtd.n5 gnd 0.236f
C515 vtd.n6 gnd 0.323f
C516 vtd.t25 gnd 2.08f
C517 vtd.t29 gnd 0.404f
C518 vtd.n7 gnd 1.27f
C519 vtd.t27 gnd 0.403f
C520 vtd.t28 gnd 0.401f
C521 vtd.n8 gnd 0.398f
C522 vtd.t26 gnd 0.401f
C523 vtd.n9 gnd 0.205f
C524 vtd.t24 gnd 0.401f
C525 vtd.t1 gnd 0.0205f
C526 vtd.t5 gnd 0.0115f
C527 vtd.n10 gnd 0.439f
C528 vtd.t2 gnd 0.0115f
C529 vtd.n11 gnd 0.236f
C530 vtd.t6 gnd 0.0115f
C531 vtd.n12 gnd 0.248f
C532 vtd.t3 gnd 0.0115f
C533 vtd.t0 gnd 0.0115f
C534 vtd.t4 gnd 0.0206f
C535 vtd.n13 gnd 0.4f
C536 vtd.t7 gnd 0.0115f
C537 vtd.n14 gnd 0.22f
C538 vtd.n15 gnd 0.324f
C539 vtd.n16 gnd 0.453f
C540 vtd.t11 gnd 0.024f
C541 vtd.t10 gnd 0.401f
C542 vtd.t8 gnd 0.401f
C543 vtd.t9 gnd 0.0229f
C544 vtd.t23 gnd 0.0229f
C545 vtd.t22 gnd 0.401f
C546 vtd.t20 gnd 0.401f
C547 vtd.t21 gnd 0.0229f
C548 vtd.t13 gnd 0.0229f
C549 vtd.t12 gnd 0.401f
C550 vtd.t14 gnd 0.401f
C551 vtd.t15 gnd 0.0229f
C552 vtd.t17 gnd 0.0229f
C553 vtd.t16 gnd 0.401f
C554 vtd.t18 gnd 0.401f
C555 vtd.t19 gnd 0.0239f
C556 vtd.n17 gnd 0.532f
C557 vtd.n18 gnd 0.341f
C558 vtd.n19 gnd 0.341f
C559 vtd.n20 gnd 0.626f
C560 vpwr.n0 gnd 6.98e-19
C561 vpwr.n1 gnd 5.16e-19
C562 vpwr.n2 gnd 0.00119f
C563 vpwr.t0 gnd 0.00306f
C564 vpwr.n3 gnd 0.00177f
C565 vpwr.n4 gnd 0.00195f
C566 vpwr.n5 gnd 8.2e-19
C567 vpwr.t31 gnd 0.00188f
C568 vpwr.n6 gnd 0.00234f
C569 vpwr.n7 gnd 0.00381f
C570 vpwr.n8 gnd 4.86e-19
C571 vpwr.n9 gnd 5.16e-19
C572 vpwr.n10 gnd 5.16e-19
C573 vpwr.n11 gnd 0.00119f
C574 vpwr.n12 gnd 0.0079f
C575 vpwr.n13 gnd 5.47e-19
C576 vpwr.t30 gnd 0.00144f
C577 vpwr.t3 gnd 0.00361f
C578 vpwr.n14 gnd 0.00619f
C579 vpwr.n15 gnd 0.00244f
C580 vpwr.n16 gnd 0.00179f
C581 vpwr.n17 gnd 3.49e-19
C582 vpwr.n18 gnd 3.21e-19
C583 vpwr.n19 gnd 7.17e-19
C584 vpwr.n20 gnd 0.00252f
C585 vpwr.n21 gnd 4.92e-19
C586 vpwr.n22 gnd 0.00241f
C587 vpwr.n23 gnd 5.75e-19
C588 vpwr.n24 gnd 6.85e-19
C589 vpwr.n25 gnd 0.00178f
C590 vpwr.n26 gnd 0.0373f
C591 vpwr.n27 gnd 0.0589f
C592 vpwr.n28 gnd 0.392f
C593 vpwr.n29 gnd 0.0742f
C594 vpwr.n30 gnd 0.00822f
C595 vpwr.t14 gnd 0.00142f
C596 vpwr.t7 gnd 0.00142f
C597 vpwr.n31 gnd 0.00306f
C598 vpwr.t27 gnd 0.00329f
C599 vpwr.n32 gnd 0.00734f
C600 vpwr.n33 gnd 0.00725f
C601 vpwr.n34 gnd 0.00151f
C602 vpwr.n35 gnd 0.00725f
C603 vpwr.n36 gnd 0.00725f
C604 vpwr.t11 gnd 0.0063f
C605 vpwr.n37 gnd 0.00257f
C606 vpwr.n38 gnd 0.00725f
C607 vpwr.t2 gnd 9.31e-19
C608 vpwr.t21 gnd 0.00176f
C609 vpwr.n39 gnd 0.00287f
C610 vpwr.n40 gnd 0.00435f
C611 vpwr.t19 gnd 0.00211f
C612 vpwr.t29 gnd 9.49e-19
C613 vpwr.n41 gnd 0.00829f
C614 vpwr.n42 gnd 0.0497f
C615 vpwr.t23 gnd 0.00277f
C616 vpwr.t9 gnd 1e-18
C617 vpwr.n43 gnd 0.00369f
C618 vpwr.n44 gnd 0.00654f
C619 vpwr.n45 gnd 0.0052f
C620 vpwr.n46 gnd 0.00352f
C621 vpwr.n47 gnd 0.0106f
C622 vpwr.n48 gnd 0.00725f
C623 vpwr.n49 gnd 0.002f
C624 vpwr.n50 gnd 0.00686f
C625 vpwr.n51 gnd 0.00204f
C626 vpwr.n52 gnd 0.00725f
C627 vpwr.n53 gnd 0.00725f
C628 vpwr.n54 gnd 0.00725f
C629 vpwr.n55 gnd 0.00247f
C630 vpwr.n56 gnd 0.0101f
C631 vpwr.n57 gnd 0.00163f
C632 vpwr.t5 gnd 9.31e-19
C633 vpwr.t17 gnd 0.00138f
C634 vpwr.n58 gnd 0.00248f
C635 vpwr.n59 gnd 0.00669f
C636 vpwr.n60 gnd 0.00142f
C637 vpwr.n61 gnd 0.00725f
C638 vpwr.n62 gnd 0.00725f
C639 vpwr.n63 gnd 0.00725f
C640 vpwr.n64 gnd 0.00257f
C641 vpwr.n65 gnd 0.00257f
C642 vpwr.n66 gnd 0.00248f
C643 vpwr.n67 gnd 0.00725f
C644 vpwr.n68 gnd 0.00725f
C645 vpwr.n69 gnd 0.00725f
C646 vpwr.n70 gnd 0.00195f
C647 vpwr.n71 gnd 0.00213f
C648 vpwr.n72 gnd 0.00905f
C649 vpwr.n73 gnd 0.00654f
C650 vpwr.n74 gnd 0.00643f
C651 vpwr.n75 gnd 0.00624f
C652 vpwr.t28 gnd 0.0505f
C653 vpwr.t18 gnd 0.0416f
C654 vpwr.t22 gnd 0.0505f
C655 vpwr.t8 gnd 0.0327f
C656 vpwr.t1 gnd 0.0253f
C657 vpwr.t20 gnd 0.0253f
C658 vpwr.t25 gnd 0.0224f
C659 vpwr.t15 gnd 0.0244f
C660 vpwr.t10 gnd 0.039f
C661 vpwr.t4 gnd 0.0387f
C662 vpwr.t16 gnd 0.0312f
C663 vpwr.t12 gnd 0.0315f
C664 vpwr.t24 gnd 0.0252f
C665 vpwr.t26 gnd 0.0473f
C666 vpwr.t13 gnd 0.0463f
C667 vpwr.t6 gnd 0.0203f
C668 vpwr.n76 gnd 0.00221f
C669 vpwr.n77 gnd 0.0549f
C670 vpwr.n78 gnd 0.00292f
C671 vpwr.n79 gnd 0.00111f
C672 vpwr.n80 gnd 0.00502f
C673 vpwr.n81 gnd 0.00164f
C674 vpwr.n82 gnd 0.00519f
C675 vpwr.n83 gnd 0.0339f
C676 sensor_0.a.n0 gnd 0.396f
C677 sensor_0.a.n1 gnd 0.413f
C678 sensor_0.a.t15 gnd 0.277f
C679 sensor_0.a.t14 gnd 0.276f
C680 sensor_0.a.n2 gnd 0.293f
C681 sensor_0.a.t12 gnd 0.276f
C682 sensor_0.a.n3 gnd 0.15f
C683 sensor_0.a.t13 gnd 0.276f
C684 sensor_0.a.n4 gnd 0.148f
C685 sensor_0.a.t1 gnd 0.0159f
C686 sensor_0.a.t0 gnd 0.276f
C687 sensor_0.a.t2 gnd 0.276f
C688 sensor_0.a.t3 gnd 0.0177f
C689 sensor_0.a.t11 gnd 0.0141f
C690 sensor_0.a.t8 gnd 0.00791f
C691 sensor_0.a.n5 gnd 0.277f
C692 sensor_0.a.t7 gnd 0.00792f
C693 sensor_0.a.n6 gnd 0.152f
C694 sensor_0.a.t4 gnd 0.00792f
C695 sensor_0.a.n7 gnd 0.19f
C696 sensor_0.a.t6 gnd 0.0141f
C697 sensor_0.a.t10 gnd 0.00791f
C698 sensor_0.a.n8 gnd 0.276f
C699 sensor_0.a.t5 gnd 0.0079f
C700 sensor_0.a.n9 gnd 0.154f
C701 sensor_0.a.t9 gnd 0.00792f
C702 sensor_0.a.n10 gnd 0.19f
C703 sensor_0.a.n11 gnd 0.384f
C704 sensor_0.b.t17 gnd 0.0077f
C705 sensor_0.b.t0 gnd 0.0077f
C706 sensor_0.b.n0 gnd 0.0683f
C707 sensor_0.b.t18 gnd 0.0077f
C708 sensor_0.b.t19 gnd 0.0077f
C709 sensor_0.b.n1 gnd 0.0506f
C710 sensor_0.b.n2 gnd 0.162f
C711 sensor_0.b.t4 gnd 0.00651f
C712 sensor_0.b.t12 gnd 0.00386f
C713 sensor_0.b.n3 gnd 0.139f
C714 sensor_0.b.t6 gnd 0.00385f
C715 sensor_0.b.n4 gnd 0.0928f
C716 sensor_0.b.t14 gnd 0.00385f
C717 sensor_0.b.n5 gnd 0.137f
C718 sensor_0.b.n6 gnd 0.202f
C719 sensor_0.b.t3 gnd 0.134f
C720 sensor_0.b.t11 gnd 0.127f
C721 sensor_0.b.t5 gnd 0.127f
C722 sensor_0.b.t13 gnd 0.0845f
C723 sensor_0.b.t32 gnd 0.134f
C724 sensor_0.b.t24 gnd 0.127f
C725 sensor_0.b.t31 gnd 0.127f
C726 sensor_0.b.t23 gnd 0.0845f
C727 sensor_0.b.t26 gnd 0.134f
C728 sensor_0.b.t34 gnd 0.127f
C729 sensor_0.b.t21 gnd 0.127f
C730 sensor_0.b.t29 gnd 0.0845f
C731 sensor_0.b.t20 gnd 0.134f
C732 sensor_0.b.t27 gnd 0.127f
C733 sensor_0.b.t28 gnd 0.127f
C734 sensor_0.b.t35 gnd 0.0845f
C735 sensor_0.b.t30 gnd 0.134f
C736 sensor_0.b.t22 gnd 0.127f
C737 sensor_0.b.t33 gnd 0.127f
C738 sensor_0.b.t25 gnd 0.0856f
C739 sensor_0.b.n7 gnd 0.119f
C740 sensor_0.b.n8 gnd 0.0626f
C741 sensor_0.b.n9 gnd 0.0626f
C742 sensor_0.b.n10 gnd 0.0626f
C743 sensor_0.b.t1 gnd 0.134f
C744 sensor_0.b.t9 gnd 0.127f
C745 sensor_0.b.t7 gnd 0.127f
C746 sensor_0.b.t15 gnd 0.0845f
C747 sensor_0.b.n11 gnd 0.0519f
C748 sensor_0.b.t2 gnd 0.00705f
C749 sensor_0.b.t10 gnd 0.00386f
C750 sensor_0.b.n12 gnd 0.138f
C751 sensor_0.b.t8 gnd 0.00386f
C752 sensor_0.b.n13 gnd 0.073f
C753 sensor_0.b.t16 gnd 0.00389f
C754 sensor_0.b.n14 gnd 0.0704f
C755 sensor_0.b.n15 gnd 0.0509f
C756 vd.t84 gnd 21.7f
C757 vd.t85 gnd 21.7f
C758 vd.t83 gnd 43.1f
C759 vd.n0 gnd 21.5f
C760 vd.n1 gnd 13.7f
C761 vd.t80 gnd 0.0573f
C762 vd.n2 gnd 17.5f
C763 vd.t23 gnd 0.00529f
C764 vd.t30 gnd 0.00264f
C765 vd.n3 gnd 0.00881f
C766 vd.t21 gnd 0.0301f
C767 vd.n4 gnd 0.191f
C768 vd.t44 gnd 0.00264f
C769 vd.t1 gnd 0.00264f
C770 vd.n5 gnd 0.0408f
C771 vd.n6 gnd 0.0645f
C772 vd.t3 gnd 0.00264f
C773 vd.t38 gnd 0.00264f
C774 vd.n7 gnd 0.0408f
C775 vd.n8 gnd 0.0539f
C776 vd.t34 gnd 0.00363f
C777 vd.n9 gnd 0.0826f
C778 vd.t72 gnd 0.00363f
C779 vd.n10 gnd 0.0782f
C780 vd.t77 gnd 0.00264f
C781 vd.t32 gnd 0.00264f
C782 vd.n11 gnd 0.0408f
C783 vd.n12 gnd 0.0488f
C784 vd.t26 gnd 0.00264f
C785 vd.t28 gnd 0.00264f
C786 vd.n13 gnd 0.0408f
C787 vd.n14 gnd 0.0445f
C788 vd.t58 gnd 0.00363f
C789 vd.n15 gnd 0.0869f
C790 vd.t56 gnd 0.00264f
C791 vd.t54 gnd 0.00264f
C792 vd.n16 gnd 0.0438f
C793 vd.n17 gnd 0.0486f
C794 vd.t52 gnd 0.00264f
C795 vd.t64 gnd 0.00264f
C796 vd.n18 gnd 0.0408f
C797 vd.n19 gnd 0.0539f
C798 vd.t62 gnd 0.00367f
C799 vd.n20 gnd 0.0913f
C800 vd.t60 gnd 0.00264f
C801 vd.t68 gnd 0.00264f
C802 vd.n21 gnd 0.0408f
C803 vd.n22 gnd 0.0437f
C804 vd.t50 gnd 0.00264f
C805 vd.t66 gnd 0.00264f
C806 vd.n23 gnd 0.0408f
C807 vd.n24 gnd 0.0368f
C808 vd.t16 gnd 0.00265f
C809 vd.t13 gnd 0.0301f
C810 vd.t48 gnd 0.00264f
C811 vd.t15 gnd 0.00264f
C812 vd.n25 gnd 0.00698f
C813 vd.n26 gnd 0.184f
C814 vd.t0 gnd 0.161f
C815 vd.t43 gnd 0.161f
C816 vd.t29 gnd 0.161f
C817 vd.t22 gnd 0.161f
C818 vd.n27 gnd 0.227f
C819 vd.n28 gnd 0.113f
C820 vd.t2 gnd 0.161f
C821 vd.t37 gnd 0.199f
C822 vd.t33 gnd 0.24f
C823 vd.t71 gnd 0.202f
C824 vd.t76 gnd 0.161f
C825 vd.t31 gnd 0.161f
C826 vd.t25 gnd 0.113f
C827 vd.n29 gnd 0.0806f
C828 vd.n30 gnd 0.0589f
C829 vd.n31 gnd 0.0589f
C830 vd.t27 gnd 0.106f
C831 vd.n32 gnd 0.118f
C832 vd.n33 gnd 0.118f
C833 vd.t51 gnd 0.161f
C834 vd.t53 gnd 0.161f
C835 vd.t55 gnd 0.161f
C836 vd.t57 gnd 0.144f
C837 vd.n34 gnd 0.121f
C838 vd.n35 gnd 0.0497f
C839 vd.n36 gnd 0.0493f
C840 vd.t63 gnd 0.199f
C841 vd.t61 gnd 0.234f
C842 vd.t59 gnd 0.196f
C843 vd.t67 gnd 0.161f
C844 vd.t49 gnd 0.161f
C845 vd.t65 gnd 0.115f
C846 vd.t47 gnd 0.106f
C847 vd.n37 gnd 0.0806f
C848 vd.n38 gnd 0.0497f
C849 vd.n39 gnd 0.181f
C850 vd.n40 gnd 0.0688f
C851 vd.t14 gnd 0.1f
C852 vd.n41 gnd 0.0806f
C853 vd.n42 gnd 0.0147f
C854 vd.n43 gnd 0.0144f
C855 vd.n44 gnd 0.0532f
C856 vd.n45 gnd 0.0143f
C857 vd.n46 gnd 0.102f
C858 vd.n47 gnd 0.0142f
C859 vd.n48 gnd 0.00352f
C860 vd.n49 gnd 0.0108f
C861 vd.n50 gnd 6.74e-19
C862 vd.t82 gnd 0.00793f
C863 vd.n51 gnd 0.00188f
C864 vd.n52 gnd 0.0124f
C865 vd.n53 gnd 0.00255f
C866 vd.n54 gnd 0.0143f
C867 vd.n55 gnd 7.28e-19
C868 vd.n56 gnd 0.00522f
C869 vd.n57 gnd 0.0143f
C870 vd.t81 gnd 0.149f
C871 vd.n59 gnd 0.0142f
C872 vd.n60 gnd 0.00522f
C873 vd.n62 gnd 0.144f
C874 vd.n63 gnd 0.0191f
C875 vd.n64 gnd 0.0142f
C876 vd.n65 gnd 0.00581f
C877 vd.n66 gnd 0.0096f
C878 vd.n67 gnd 0.125f
C879 vd.n68 gnd 0.0097f
C880 vd.n69 gnd 0.00593f
C881 vd.n70 gnd 0.0151f
C882 vd.n71 gnd 0.0302f
C883 vd.n72 gnd 0.0153f
C884 vd.n73 gnd 0.00837f
C885 vd.n74 gnd 0.0461f
C886 vd.n75 gnd 0.00327f
C887 vd.n76 gnd 0.00883f
C888 vd.n77 gnd 0.00182f
C889 vd.n78 gnd 0.00237f
C890 vd.n79 gnd 0.00219f
C891 vd.n80 gnd 0.0106f
C892 vd.n81 gnd 0.014f
C893 vd.n82 gnd 0.135f
C894 vd.t19 gnd 0.00556f
C895 vd.t20 gnd 0.00552f
C896 vd.t70 gnd 0.0058f
C897 vd.n83 gnd 0.0893f
C898 vd.t17 gnd 0.0924f
C899 vd.n84 gnd 0.0732f
C900 vd.n85 gnd 0.109f
C901 vd.n86 gnd 0.0576f
C902 vd.n87 gnd 0.291f
C903 vd.n88 gnd 0.232f
C904 vd.n89 gnd 0.019f
C905 vd.n90 gnd 0.019f
C906 vd.t42 gnd 0.0941f
C907 vd.t18 gnd 0.102f
C908 vd.t35 gnd 0.349f
C909 vd.n91 gnd 0.278f
C910 vd.n92 gnd 0.0108f
C911 vd.t4 gnd 0.156f
C912 vd.n93 gnd 0.196f
C913 vd.n94 gnd 0.0142f
C914 vd.n95 gnd 0.014f
C915 vd.n96 gnd 0.0119f
C916 vd.t12 gnd 0.00558f
C917 vd.t9 gnd 0.0924f
C918 vd.t11 gnd 0.00563f
C919 vd.t46 gnd 0.00588f
C920 vd.n97 gnd 0.102f
C921 vd.n98 gnd 0.0671f
C922 vd.n99 gnd 0.0801f
C923 vd.n100 gnd 0.00177f
C924 vd.t8 gnd 0.00529f
C925 vd.n101 gnd 0.0307f
C926 vd.t7 gnd 0.00556f
C927 vd.t74 gnd 0.00528f
C928 vd.t41 gnd 0.00528f
C929 vd.n102 gnd 0.0419f
C930 vd.n103 gnd 0.0544f
C931 vd.t5 gnd 0.0924f
C932 vd.n104 gnd 0.0612f
C933 vd.n105 gnd 0.00621f
C934 vd.n106 gnd 0.00285f
C935 vd.n107 gnd 0.051f
C936 vd.n108 gnd 0.0593f
C937 vd.n109 gnd 0.348f
C938 vd.t6 gnd 0.236f
C939 vd.n110 gnd 0.288f
C940 vd.n111 gnd 0.0224f
C941 vd.n112 gnd 0.0223f
C942 vd.t73 gnd 0.425f
C943 vd.t40 gnd 0.265f
C944 vd.n113 gnd 0.196f
C945 vd.n114 gnd 0.0141f
C946 vd.n115 gnd 0.0152f
C947 vd.n116 gnd 0.119f
C948 vd.n117 gnd 0.142f
C949 vd.t24 gnd 0.103f
C950 vd.t45 gnd 0.0819f
C951 vd.n118 gnd 0.0846f
C952 vd.n119 gnd 0.0846f
C953 vd.n120 gnd 0.17f
C954 vd.n121 gnd 0.00604f
C955 vd.n122 gnd 0.00602f
C956 vd.t78 gnd 0.252f
C957 vd.n123 gnd 0.29f
C958 vd.n124 gnd 0.0173f
C959 vd.n125 gnd 0.0171f
C960 vd.t79 gnd 0.137f
C961 vd.t75 gnd 0.273f
C962 vd.t10 gnd 0.173f
C963 vd.n126 gnd 0.118f
C964 vd.n127 gnd 0.0115f
C965 vd.n128 gnd 0.0125f
C966 vd.n129 gnd 0.117f
C967 vd.n130 gnd 0.293f
C968 vd.n131 gnd 0.00929f
C969 vd.n132 gnd 0.00918f
C970 vd.t69 gnd 0.196f
C971 vd.t36 gnd 0.193f
C972 vd.t39 gnd 0.296f
C973 vd.n133 gnd 0.196f
C974 vd.n134 gnd 0.0132f
C975 vd.n135 gnd 0.0143f
C976 vd.n136 gnd 0.166f
C977 vd.n137 gnd 0.0961f
C978 vd.n138 gnd 0.563f
C979 vd.n139 gnd 1.81f
C980 vd.n140 gnd 5.37f
C981 vd.n141 gnd 4.9f
C982 vd.n142 gnd 0.461f
C983 buffer_0.a.n0 gnd 1.52f
C984 buffer_0.a.n1 gnd 1.5f
C985 buffer_0.a.t11 gnd 0.0207f
C986 buffer_0.a.t21 gnd 0.514f
C987 buffer_0.a.t22 gnd 0.509f
C988 buffer_0.a.n2 gnd 0.575f
C989 buffer_0.a.t23 gnd 0.509f
C990 buffer_0.a.n3 gnd 0.295f
C991 buffer_0.a.t24 gnd 0.509f
C992 buffer_0.a.n4 gnd 0.295f
C993 buffer_0.a.t19 gnd 0.509f
C994 buffer_0.a.n5 gnd 0.295f
C995 buffer_0.a.t10 gnd 0.509f
C996 buffer_0.a.t20 gnd 0.509f
C997 buffer_0.a.t17 gnd 0.509f
C998 buffer_0.a.t25 gnd 0.509f
C999 buffer_0.a.t18 gnd 0.509f
C1000 buffer_0.a.t26 gnd 0.514f
C1001 buffer_0.a.n6 gnd 0.574f
C1002 buffer_0.a.n7 gnd 0.295f
C1003 buffer_0.a.n8 gnd 0.295f
C1004 buffer_0.a.n9 gnd 0.311f
C1005 buffer_0.a.n10 gnd 0.291f
C1006 buffer_0.a.n11 gnd 0.0789f
C1007 buffer_0.a.n12 gnd 0.352f
C1008 buffer_0.a.t12 gnd 0.393f
C1009 buffer_0.a.t13 gnd 0.0421f
C1010 buffer_0.a.t5 gnd 0.0207f
C1011 buffer_0.a.t8 gnd 0.0207f
C1012 buffer_0.a.t4 gnd 0.0207f
C1013 buffer_0.a.n13 gnd 0.304f
C1014 buffer_0.a.n14 gnd 0.582f
C1015 buffer_0.a.t0 gnd 0.0207f
C1016 buffer_0.a.t6 gnd 0.0207f
C1017 buffer_0.a.n15 gnd 0.302f
C1018 buffer_0.a.n16 gnd 0.515f
C1019 buffer_0.a.t9 gnd 0.0207f
C1020 buffer_0.a.t3 gnd 0.0207f
C1021 buffer_0.a.n17 gnd 0.304f
C1022 buffer_0.a.n18 gnd 0.384f
C1023 buffer_0.a.t7 gnd 0.0207f
C1024 buffer_0.a.t2 gnd 0.0207f
C1025 buffer_0.a.n19 gnd 0.301f
C1026 buffer_0.a.t14 gnd 0.398f
C1027 buffer_0.a.t1 gnd 0.0207f
C1028 buffer_0.a.t15 gnd 0.0207f
C1029 buffer_0.a.t16 gnd 0.0207f
C1030 buffer_0.a.n20 gnd 0.486f
C1031 buffer_0.a.n21 gnd 0.293f
C1032 out_buff.t4 gnd 0.00405f
C1033 out_buff.t10 gnd 0.00405f
C1034 out_buff.n0 gnd 0.0553f
C1035 out_buff.t14 gnd 0.00405f
C1036 out_buff.t17 gnd 0.00405f
C1037 out_buff.n1 gnd 0.0913f
C1038 out_buff.t0 gnd 0.00405f
C1039 out_buff.t1 gnd 0.00405f
C1040 out_buff.n2 gnd 0.0627f
C1041 out_buff.n3 gnd 0.0812f
C1042 out_buff.t16 gnd 0.00557f
C1043 out_buff.n4 gnd 0.126f
C1044 out_buff.t18 gnd 0.00405f
C1045 out_buff.t20 gnd 0.00405f
C1046 out_buff.n5 gnd 0.0627f
C1047 out_buff.t15 gnd 0.00405f
C1048 out_buff.t12 gnd 0.00405f
C1049 out_buff.n6 gnd 0.0672f
C1050 out_buff.t13 gnd 0.00949f
C1051 out_buff.n7 gnd 0.174f
C1052 out_buff.n8 gnd 0.0565f
C1053 out_buff.n9 gnd 0.084f
C1054 out_buff.t5 gnd 0.00405f
C1055 out_buff.t2 gnd 0.00405f
C1056 out_buff.n10 gnd 0.0599f
C1057 out_buff.t6 gnd 0.00405f
C1058 out_buff.t9 gnd 0.00405f
C1059 out_buff.n11 gnd 0.0553f
C1060 out_buff.t8 gnd 0.00405f
C1061 out_buff.t11 gnd 0.00405f
C1062 out_buff.n12 gnd 0.0545f
C1063 out_buff.t7 gnd 0.00405f
C1064 out_buff.t3 gnd 0.00405f
C1065 out_buff.n13 gnd 0.104f
C1066 out_buff.n14 gnd 0.115f
C1067 out_buff.n15 gnd 0.101f
C1068 out_buff.n16 gnd 0.0653f
C1069 out_buff.n17 gnd 0.0964f
C1070 out_buff.n18 gnd 0.0578f
C1071 out_buff.t28 gnd 50.3f
C1072 out_buff.n19 gnd 0.211f
C1073 out_buff.t25 gnd 0.0766f
C1074 out_buff.t24 gnd 0.0833f
C1075 out_buff.t23 gnd 0.077f
C1076 out_buff.n20 gnd 0.151f
C1077 out_buff.t30 gnd 0.0783f
C1078 out_buff.n21 gnd 0.0777f
C1079 out_buff.t29 gnd 0.0776f
C1080 out_buff.n22 gnd 0.079f
C1081 out_buff.t21 gnd 0.0773f
C1082 out_buff.n23 gnd 0.0785f
C1083 out_buff.t26 gnd 0.076f
C1084 out_buff.n24 gnd 0.0815f
C1085 out_buff.t27 gnd 0.0765f
C1086 out_buff.n25 gnd 0.0807f
C1087 out_buff.t31 gnd 0.078f
C1088 out_buff.n26 gnd 0.0785f
C1089 out_buff.t22 gnd 0.0778f
C1090 out_buff.n27 gnd 0.0783f
C1091 out_buff.n28 gnd 0.118f
C1092 out_buff.n29 gnd 0.142f
C1093 out_buff.t19 gnd 0.0847f
C1094 out_buff.n30 gnd 0.337f
C1095 out_buff.n31 gnd 1.14f
.ends

