magic
tech sky130A
timestamp 1644072167
<< metal4 >>
rect 4400 4400 8600 4900
<< metal5 >>
rect 0 7600 8100 8100
rect 0 6800 7300 7300
rect 0 500 500 6800
rect 800 6000 6500 6500
rect 800 1300 1300 6000
rect 1600 5200 5700 5700
rect 1600 2100 2100 5200
rect 2400 4400 4900 4900
rect 2400 2900 2900 4400
rect 5200 2900 5700 5200
rect 2400 2400 5700 2900
rect 6000 2100 6500 6000
rect 1600 1600 6500 2100
rect 6800 1300 7300 6800
rect 800 800 7300 1300
rect 7600 500 8100 7600
rect 0 0 8100 500
<< labels >>
flabel metal5 229 7860 229 7860 0 FreeSans 800 0 0 0 p1
port 0 nsew
flabel metal4 8326 4641 8343 4641 0 FreeSans 800 0 0 0 p2
port 2 nsew
<< end >>
