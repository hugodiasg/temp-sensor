magic
tech sky130A
magscale 1 2
timestamp 1675896714
<< metal4 >>
rect 50330 53014 53018 53018
rect 50330 52912 62561 53014
rect 50330 50436 50436 52912
rect 52912 50436 62561 52912
rect 50330 50334 62561 50436
rect 50330 50330 53018 50334
<< via4 >>
rect 50436 50436 52912 52912
<< metal5 >>
rect 56514 59194 59194 59200
rect 42526 56514 59194 59194
rect 43204 56104 45884 56109
rect 53424 56104 56104 56110
rect 43199 53424 56109 56104
rect 43204 45884 45884 53424
rect 46294 53014 48974 53018
rect 50330 53014 53018 53018
rect 46290 52912 53018 53014
rect 46290 50436 50436 52912
rect 52912 50436 53018 52912
rect 46290 50334 53018 50436
rect 46294 48974 48974 50334
rect 50330 50330 53018 50334
rect 53424 48974 56104 53424
rect 46290 46294 56110 48974
rect 46294 46290 48974 46294
rect 53424 46290 56104 46294
rect 56514 45884 59194 56514
rect 43200 43204 59200 45884
rect 43204 43199 45884 43204
rect 56514 43200 59194 43204
<< end >>
