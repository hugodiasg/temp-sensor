magic
tech sky130A
magscale 1 2
timestamp 1644599756
<< metal4 >>
rect -2499 7319 2499 7360
rect -2499 2561 2243 7319
rect 2479 2561 2499 7319
rect -2499 2520 2499 2561
rect -2499 2379 2499 2420
rect -2499 -2379 2243 2379
rect 2479 -2379 2499 2379
rect -2499 -2420 2499 -2379
rect -2499 -2561 2499 -2520
rect -2499 -7319 2243 -2561
rect 2479 -7319 2499 -2561
rect -2499 -7360 2499 -7319
<< via4 >>
rect 2243 2561 2479 7319
rect 2243 -2379 2479 2379
rect 2243 -7319 2479 -2561
<< mimcap2 >>
rect -2399 7220 2241 7260
rect -2399 2660 -1903 7220
rect 1745 2660 2241 7220
rect -2399 2620 2241 2660
rect -2399 2280 2241 2320
rect -2399 -2280 -1903 2280
rect 1745 -2280 2241 2280
rect -2399 -2320 2241 -2280
rect -2399 -2660 2241 -2620
rect -2399 -7220 -1903 -2660
rect 1745 -7220 2241 -2660
rect -2399 -7260 2241 -7220
<< mimcap2contact >>
rect -1903 2660 1745 7220
rect -1903 -2280 1745 2280
rect -1903 -7220 1745 -2660
<< metal5 >>
rect -239 7244 81 7410
rect 2201 7319 2521 7410
rect -1927 7220 1769 7244
rect -1927 2660 -1903 7220
rect 1745 2660 1769 7220
rect -1927 2636 1769 2660
rect -239 2304 81 2636
rect 2201 2561 2243 7319
rect 2479 2561 2521 7319
rect 2201 2379 2521 2561
rect -1927 2280 1769 2304
rect -1927 -2280 -1903 2280
rect 1745 -2280 1769 2280
rect -1927 -2304 1769 -2280
rect -239 -2636 81 -2304
rect 2201 -2379 2243 2379
rect 2479 -2379 2521 2379
rect 2201 -2561 2521 -2379
rect -1927 -2660 1769 -2636
rect -1927 -7220 -1903 -2660
rect 1745 -7220 1769 -2660
rect -1927 -7244 1769 -7220
rect -239 -7410 81 -7244
rect 2201 -7319 2243 -2561
rect 2479 -7319 2521 -2561
rect 2201 -7410 2521 -7319
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2499 2520 2341 7360
string parameters w 23.2 l 23.2 val 1.094k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
