** sch_path: /foss/designs/temp-sensor/device-complete/xschem/device-complete-tb.sch
**.subckt device-complete-tb
vpwr vpwr GND 1.8
V3 clk GND pulse 0 1.8 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 '
vdd vd GND 1.8
ibias vd ib 1u
VSS vs GND 0
x1 vd clk out vpwr ib net1 GND device-complete-pex
**** begin user architecture code

*cmd step stop

.save
.control
destroy all
save all
set color0=white
set color1=black
set temp=60
set hcopypscolor = 1
set wr_singlescale
option numdgt=7
tran 40p 10u
*let pot=-i(vdd)*vd
save all

plot x1.vts x1.out_sigma x1.out_buf
*plot x1.vts x1.out_buf
plot out


*meas tran pot_avg avg pot from=0 to=5u
*plot pot pot_avg pot_rms

*wrdata ./tran10.txt x1.vts x1.out_sigma out

*linearize out
*fft out
*hardcopy ~/fft56.ps mag(out_ask) xlimit 1G 4G ylimit 0 55u
*plot mag(out) xlimit 1G 4G ylimit 0 65u

*wrdata ./fft10.txt mag(out)




.endc



 .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/temp-sensor/device-complete/xschem/device-complete-pex.sym # of
*+ pins=7
** sym_path: /foss/designs/temp-sensor/device-complete/xschem/device-complete-pex.sym
** sch_path: /foss/designs/temp-sensor/device-complete/xschem/device-complete-pex.sch
.subckt device-complete-pex vd clk out vpwr ib ib2 gnd
*.iopin vd
*.ipin clk
*.opin out
*.iopin vpwr
*.iopin ib
*.iopin ib2
*.iopin gnd
**** begin user architecture code



* NGSPICE file created from device-complete.ext - technology: sky130A

*.subckt device-complete gnd clk ib vd out vpwr
X0 gnd.t77 buffer_0.d out_buff.t2 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X1 a_16688_5320# a_16854_3988# gnd.t82 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X2 vd.t22 buffer_0.a.t17 buffer_0.d vd.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X3 sensor_0.a.t11 sensor_0.b.t20 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X4 out_buff.t4 buffer_0.d gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X5 sensor_0.b.t17 sensor_0.b.t16 gnd.t89 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X6 a_15868_2881# a_14791_2515# a_15706_2515# vpwr.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69
+ as=0.0588 ps=0.7 w=0.42 l=0.15
X7 gnd.t137 vpwr.t30 a_15403_2515# gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441
+ ps=0.63 w=0.42 l=0.15
X8 a_15546_5320# a_15712_3988# gnd.t8 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X9 vd.t20 buffer_0.a.t18 buffer_0.d vd.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X10 buffer_0.a.t4 buffer_0.a.t2 buffer_0.a.t3 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0
+ ps=0 w=1 l=1
X11 gnd.t14 sensor_0.b.t21 vtd.t23 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X12 a_15141_2515# a_14791_2515# a_15046_2515# vpwr.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0724
+ pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X13 sensor_0.c sensor_0.c sensor_0.c vd.t80 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6
+ w=2 l=1
X14 buffer_0.c.t9 vts.t25 buffer_0.b.t8 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X15 gnd.t171 gnd.t169 gnd.t170 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X16 a_14550_5320# a_14716_3988# gnd.t30 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X17 a_15815_2515# a_14625_2515# a_15706_2515# gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75
+ as=0.0711 ps=0.755 w=0.36 l=0.15
X18 vd.t18 buffer_0.a.t19 buffer_0.d vd.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58
+ w=1 l=1
X19 buffer_0.c.t19 out_buff.t21 buffer_0.a.t16 gnd.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X20 gnd.t33 sensor_0.b.t14 sensor_0.b.t15 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X21 vts.t24 vtd.t12 vtd.t13 vts.t23 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X22 a_16356_5320# a_16522_3988# gnd.t7 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X23 vd.t55 vd.t53 vd.t55 vd.t54 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X24 buffer_0.c.t8 vts.t26 buffer_0.b.t2 gnd.t36 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X25 gnd.t10 ib.t3 ib.t4 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 buffer_0.d buffer_0.d gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X27 gnd.t168 gnd.t166 gnd.t167 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X28 vtd.t11 vtd.t10 vts.t22 vts.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 gnd.t115 sensor_0.b.t22 sensor_0.a.t10 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X30 vd.t78 buffer_0.b.t10 out_buff.t20 vd.t77 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X31 gnd.t165 gnd.t163 gnd.t164 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X32 vtd.t22 sensor_0.b.t23 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1
+ l=1
X33 out_sigma.t0 a_16445_2515# vpwr.t11 vpwr.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52
+ as=0.154 ps=1.34 w=1 l=0.15
X34 gnd.t71 buffer_0.d out_buff.t1 gnd.t70 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X35 vts.t20 vtd.t14 vtd.t15 vts.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 buffer_0.c.t18 out_buff.t22 buffer_0.a.t15 gnd.t105 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X37 vtd.t21 sensor_0.b.t24 gnd.t109 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X38 vpwr.t23 clk.t0 a_14625_2515# vpwr.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166
+ ps=1.8 w=0.64 l=0.15
X39 out_buff.t5 buffer_0.d gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X40 a_17020_5320# sigma-delta_0.x1.Q gnd.t129 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X41 a_15237_2515# a_14791_2515# a_15141_2515# gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1
+ as=0.0594 ps=0.69 w=0.36 l=0.15
X42 a_15706_2515# a_14625_2515# a_15359_2757# vpwr.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7
+ as=0.129 ps=1.18 w=0.42 l=0.15
X43 vtd.t7 vtd.t6 vts.t18 vts.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X44 vd.t0 a_6126_29386# gnd.t24 sky130_fd_pr__res_xhigh_po_0p35 l=5
X45 sensor_0.b.t18 vtd.t24 sensor_0.c vd.t79 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58
+ w=2 l=1
X46 a_15359_2757# a_15141_2515# vpwr.t21 vpwr.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18
+ as=0.218 ps=2.2 w=0.84 l=0.15
X47 gnd.t35 clk.t1 a_14625_2515# gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36
+ w=0.42 l=0.15
X48 buffer_0.a.t6 buffer_0.a.t5 vd.t16 vd.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X49 gnd.t12 sensor_0.b.t12 sensor_0.b.t13 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X50 vpwr.t19 a_15706_2515# a_15881_2489# vpwr.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67
+ as=0.0567 ps=0.69 w=0.42 l=0.15
X51 vts.t16 vtd.t8 vtd.t9 vts.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X52 a_15046_2515# sigma-delta_0.x1.D vpwr.t13 vpwr.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73
+ as=0.109 ps=1.36 w=0.42 l=0.15
X53 vd.t35 sensor_0.a.t2 sensor_0.a.t3 vd.t34 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58
+ ps=4.58 w=2 l=1
X54 gnd.t67 buffer_0.d buffer_0.d gnd.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X55 a_15881_2489# a_15706_2515# a_16060_2515# gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36
+ as=0.064 ps=0.725 w=0.42 l=0.15
X56 buffer_0.a.t8 out_buff.t23 buffer_0.c.t17 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X57 sensor_0.b.t11 sensor_0.b.t10 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X58 a_14882_5320# a_15048_3988# gnd.t78 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X59 buffer_0.d buffer_0.a.t20 vd.t14 vd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29
+ w=1 l=1
X60 gnd.t140 sensor_0.b.t25 sensor_0.a.t9 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X61 buffer_0.c.t7 vts.t27 buffer_0.b.t3 gnd.t135 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X62 buffer_0.c.t6 vts.t28 buffer_0.b.t6 gnd.t138 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X63 buffer_0.b.t7 vts.t29 buffer_0.c.t5 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X64 buffer_0.b.t0 vts.t30 buffer_0.c.t4 gnd.t120 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X65 sigma-delta_0.x1.Q a_15881_2489# gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82
+ as=0.169 ps=1.82 w=0.65 l=0.15
X66 vd.t12 buffer_0.a.t21 buffer_0.d vd.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29
+ w=1 l=1
X67 buffer_0.c.t20 ib.t5 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29
+ w=1 l=1
X68 vts.t7 vts.t4 vts.t6 vts.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X69 buffer_0.c.t16 out_buff.t24 buffer_0.a.t9 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X70 gnd.t65 buffer_0.d buffer_0.d gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58
+ w=1 l=1
X71 gnd.t63 buffer_0.d buffer_0.d gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X72 a_15359_2757# a_15141_2515# gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135
+ ps=1.15 w=0.64 l=0.15
X73 vpwr.t17 a_15359_2757# a_15249_2881# vpwr.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755
+ as=0.116 ps=0.97 w=0.42 l=0.15
X74 buffer_0.d buffer_0.a.t22 vd.t10 vd.t9 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X75 a_15706_2515# a_14791_2515# a_15359_2757# gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755
+ as=0.0999 ps=0.985 w=0.36 l=0.15
X76 gnd.t144 sensor_0.b.t26 vtd.t20 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X77 vd.t25 vtd.t25 vts.t14 vd.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X78 vd.t8 buffer_0.a.t23 buffer_0.d vd.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X79 a_15214_5320# a_15380_3988# gnd.t27 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X80 vd.t52 vd.t49 vd.t51 vd.t50 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X81 buffer_0.d buffer_0.a.t24 vd.t6 vd.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X82 buffer_0.a.t1 buffer_0.a.t0 buffer_0.a.t1 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0
+ ps=0 w=1 l=1
X83 gnd.t162 gnd.t160 gnd.t161 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X84 sensor_0.c vtd.t26 sensor_0.b.t0 vd.t23 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29
+ w=2 l=1
X85 buffer_0.a.t13 out_buff.t25 buffer_0.c.t15 gnd.t102 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X86 out_sigma.t1 a_16445_2515# gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1
+ ps=0.985 w=0.65 l=0.15
X87 buffer_0.d buffer_0.d gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X88 sensor_0.a.t8 sensor_0.b.t27 gnd.t88 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X89 sensor_0.a.t7 sensor_0.b.t28 gnd.t114 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X90 sigma-delta_0.x1.Q a_15881_2489# vpwr.t29 vpwr.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56
+ as=0.213 ps=1.67 w=1 l=0.15
X91 sensor_0.a.t1 sensor_0.a.t0 vd.t31 vd.t30 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29
+ ps=2.29 w=2 l=1
X92 gnd.t59 buffer_0.d out_buff.t6 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X93 vd.t83 out.t3 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X94 a_16060_2515# vpwr.t31 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125
+ ps=1.01 w=0.42 l=0.15
X95 vd.t48 vd.t45 vd.t47 vd.t46 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X96 out_buff.t3 buffer_0.d gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X97 a_16024_5320# a_16190_3988# gnd.t87 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X98 sensor_0.b.t9 sensor_0.b.t8 gnd.t145 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X99 gnd.t117 sensor_0.b.t29 vtd.t19 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X100 vd.t72 buffer_0.b.t11 out_buff.t18 vd.t71 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29
+ ps=2.58 w=1 l=1
X101 a_16688_5320# a_16522_3988# gnd.t26 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X102 vd.t44 vd.t41 vd.t43 vd.t42 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X103 buffer_0.a.t10 out_buff.t26 buffer_0.c.t14 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X104 sensor_0.c sensor_0.a.t12 sensor_0.d vd.t26 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29
+ ps=2.29 w=2 l=1
X105 sensor_0.d sensor_0.a.t13 sensor_0.c vd.t81 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58
+ ps=4.58 w=2 l=1
X106 a_15546_5320# a_15380_3988# gnd.t17 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X107 vpwr.t27 a_15881_2489# a_15868_2881# vpwr.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81
+ as=0.0567 ps=0.69 w=0.42 l=0.15
X108 buffer_0.c.t13 out_buff.t27 buffer_0.a.t11 gnd.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X109 gnd.t159 gnd.t157 gnd.t158 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X110 gnd.t156 gnd.t154 gnd.t155 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X111 gnd.t153 gnd.t150 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X112 vd.t40 vd.t37 vd.t39 vd.t38 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X113 buffer_0.d buffer_0.d gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X114 a_15046_2515# sigma-delta_0.x1.D gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745
+ as=0.221 ps=1.89 w=0.42 l=0.15
X115 gnd.t141 sensor_0.b.t6 sensor_0.b.t7 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X116 vtd.t1 vtd.t0 vts.t13 vts.t12 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X117 vd.t76 buffer_0.b.t12 out_buff.t19 vd.t75 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29
+ ps=2.58 w=1 l=1
X118 gnd.t53 buffer_0.d out_buff.t7 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X119 gnd.t51 buffer_0.d out_buff.t9 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X120 gnd.t139 sensor_0.b.t30 sensor_0.a.t6 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X121 a_15141_2515# a_14625_2515# a_15046_2515# gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69
+ as=0.066 ps=0.745 w=0.36 l=0.15
X122 vts.t11 vtd.t4 vtd.t5 vts.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X123 vtd.t18 sensor_0.b.t31 gnd.t142 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X124 buffer_0.b buffer_0.b.t9 vd.t74 vd.t73 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X125 out_buff.t8 buffer_0.d gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X126 out_buff.t28 buffer_0.d sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X127 a_16356_5320# a_16190_3988# gnd.t113 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X128 out_buff.t10 buffer_0.d gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X129 vtd.t3 vtd.t2 vts.t9 vts.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X130 vtd.t17 sensor_0.b.t32 gnd.t143 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X131 vd.t33 a_15712_3988# sigma-delta_0.x1.D vd.t32 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87
+ ps=6.58 w=3 l=0.15
X132 sensor_0.c vtd.t27 sensor_0.b.t19 vd.t82 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29
+ ps=2.29 w=2 l=1
X133 a_15214_5320# a_15048_3988# gnd.t131 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X134 vd.t84 out.t2 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X135 vd.t70 buffer_0.b.t13 out_buff.t17 vd.t69 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X136 buffer_0.d buffer_0.a.t25 vd.t4 vd.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X137 sensor_0.b.t1 vtd.t28 sensor_0.c vd.t36 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29
+ w=2 l=1
X138 a_17020_5320# a_16854_3988# gnd.t6 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X139 out_buff.t16 buffer_0.b.t14 vd.t68 vd.t67 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X140 gnd.t116 sensor_0.b.t4 sensor_0.b.t5 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X141 sensor_0.d vtd.t29 vd.t28 vd.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2
+ l=1
X142 buffer_0.d buffer_0.d buffer_0.d gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=2.03
+ ps=18.1 w=1 l=1
X143 a_14791_2515# a_14625_2515# vpwr.t2 vpwr.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8
+ as=0.0864 ps=0.91 w=0.64 l=0.15
X144 a_14882_5320# a_14716_3988# gnd.t95 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X145 gnd.t94 a_15712_3988# sigma-delta_0.x1.D gnd.t93 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58
+ as=0.29 ps=2.58 w=1 l=0.15
X146 sensor_0.d sensor_0.a.t14 sensor_0.c vd.t56 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29
+ ps=2.29 w=2 l=1
X147 buffer_0.a.t14 out_buff.t29 buffer_0.c.t12 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X148 buffer_0.d buffer_0.a.t26 vd.t2 vd.t1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X149 vts.t3 vts.t0 vts.t2 vts.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X150 ib.t2 ib.t0 ib.t1 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X151 a_14791_2515# a_14625_2515# gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567
+ ps=0.69 w=0.42 l=0.15
X152 a_15249_2881# a_14625_2515# a_15141_2515# vpwr.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97
+ as=0.0724 ps=0.765 w=0.42 l=0.15
X153 buffer_0.c.t3 vts.t31 buffer_0.b.t1 gnd.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X154 sensor_0.b.t3 sensor_0.b.t2 gnd.t96 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X155 gnd.t84 sensor_0.b.t33 sensor_0.a.t5 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X156 a_16024_5320# a_15712_3988# gnd.t80 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X157 out_buff.t15 buffer_0.b.t15 vd.t66 vd.t65 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X158 buffer_0.b.t4 vts.t32 buffer_0.c.t2 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X159 buffer_0.b.t5 vts.t33 buffer_0.c.t1 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X160 vd.t85 out.t1 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X161 vd.t64 buffer_0.b.t16 out_buff.t14 vd.t63 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145
+ ps=1.29 w=1 l=1
X162 gnd.t108 out_sigma.t2 out.t0 gnd.t107 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58
+ w=2 l=0.15
X163 vd.t62 buffer_0.b.t17 out_buff.t13 vd.t61 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X164 sensor_0.c sensor_0.a.t15 sensor_0.d vd.t29 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29
+ ps=2.29 w=2 l=1
X165 gnd.t134 sensor_0.b.t34 vtd.t16 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58
+ w=1 l=1
X166 out_buff.t12 buffer_0.b.t18 vd.t60 vd.t59 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X167 buffer_0.c.t11 out_buff.t30 buffer_0.a.t7 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X168 gnd.t44 buffer_0.d buffer_0.d gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X169 gnd.t42 buffer_0.d buffer_0.d gnd.t41 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X170 gnd.t126 a_15881_2489# a_15815_2515# gnd.t125 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01
+ as=0.0669 ps=0.75 w=0.42 l=0.15
X171 out_buff.t11 buffer_0.b.t19 vd.t58 vd.t57 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X172 a_15403_2515# a_15359_2757# a_15237_2515# gnd.t79 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63
+ as=0.14 ps=1.1 w=0.42 l=0.15
X173 buffer_0.d buffer_0.d gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X174 a_15249_2881# vpwr.t7 vpwr.t9 vpwr.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703
+ ps=0.755 w=0.42 l=0.15
X175 buffer_0.b.t2 vts.t34 buffer_0.c.t0 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145
+ ps=1.29 w=1 l=1
X176 a_15881_2489# vpwr.t4 vpwr.t6 vpwr.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819
+ ps=0.81 w=0.42 l=0.15
X177 a_14550_5320# out_buff.t0 gnd.t18 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X178 gnd.t124 a_15881_2489# a_16445_2515# gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109
+ ps=1.36 w=0.42 l=0.15
X179 sensor_0.a.t4 sensor_0.b.t35 gnd.t133 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29
+ ps=2.58 w=1 l=1
X180 vpwr.t25 a_15881_2489# a_16445_2515# vpwr.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34
+ as=0.166 ps=1.8 w=0.64 l=0.15
X181 buffer_0.a.t12 out_buff.t31 buffer_0.c.t10 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29
+ as=0.145 ps=1.29 w=1 l=1
X182 buffer_0.d buffer_0.d gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29
+ w=1 l=1
X183 gnd.t149 gnd.t146 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X184 a_15712_3988# gnd.t92 sky130_fd_pr__cap_mim_m3_1 l=27.2 w=27.2
R0 out_buff.n7 out_buff.t18 30.2161
R1 out_buff.n4 out_buff.t19 29.2293
R2 out_buff.n5 out_buff.t14 28.5655
R3 out_buff.n5 out_buff.t12 28.5655
R4 out_buff.n6 out_buff.t17 28.5655
R5 out_buff.n6 out_buff.t16 28.5655
R6 out_buff.n2 out_buff.t13 28.5655
R7 out_buff.n2 out_buff.t11 28.5655
R8 out_buff.n1 out_buff.t20 28.5655
R9 out_buff.n1 out_buff.t15 28.5655
R10 out_buff.n20 out_buff.t24 26.8319
R11 out_buff.n21 out_buff.t30 25.9449
R12 out_buff.n26 out_buff.t31 25.7428
R13 out_buff.n27 out_buff.t22 25.5407
R14 out_buff.n22 out_buff.t29 25.3386
R15 out_buff.n23 out_buff.t21 25.1365
R16 out_buff.n20 out_buff.t23 24.9306
R17 out_buff.n28 out_buff.t25 24.696
R18 out_buff.n25 out_buff.t27 24.5271
R19 out_buff.n24 out_buff.t26 24.1037
R20 out_buff.n0 out_buff.t6 17.4005
R21 out_buff.n0 out_buff.t3 17.4005
R22 out_buff.n10 out_buff.t2 17.4005
R23 out_buff.n10 out_buff.t4 17.4005
R24 out_buff.n11 out_buff.t9 17.4005
R25 out_buff.n11 out_buff.t10 17.4005
R26 out_buff.n12 out_buff.t1 17.4005
R27 out_buff.n12 out_buff.t5 17.4005
R28 out_buff.n13 out_buff.t7 17.4005
R29 out_buff.n13 out_buff.t8 17.4005
R30 out_buff.n30 out_buff.t0 9.50608
R31 out_buff.n14 out_buff.n13 2.74907
R32 out_buff.n17 out_buff.n9 2.41728
R33 out_buff.n24 out_buff.n23 2.30343
R34 out_buff.n22 out_buff.n21 2.29903
R35 out_buff.n28 out_buff.n27 2.2903
R36 out_buff.n26 out_buff.n25 2.25283
R37 out_buff.n16 out_buff.n15 2.1255
R38 out_buff.n15 out_buff.n14 2.1255
R39 out_buff.n29 out_buff.n19 1.97968
R40 out_buff.n18 out_buff.n17 1.83383
R41 out_buff.n3 out_buff.n1 1.74765
R42 out_buff.n19 out_buff.t28 1.69869
R43 out_buff out_buff.n29 1.51612
R44 out_buff.n30 out_buff 1.37175
R45 out_buff.n29 out_buff.n28 1.24394
R46 out_buff.n8 out_buff.n7 1.04217
R47 out_buff.n4 out_buff.n3 1.0005
R48 out_buff.n9 out_buff.n4 0.938
R49 out_buff.n25 out_buff.n24 0.680308
R50 out_buff.n23 out_buff.n22 0.678839
R51 out_buff.n27 out_buff.n26 0.678839
R52 out_buff.n8 out_buff.n5 0.664316
R53 out_buff.n3 out_buff.n2 0.664316
R54 out_buff.n9 out_buff.n8 0.646333
R55 out_buff.n21 out_buff.n20 0.63023
R56 out_buff.n7 out_buff.n6 0.610444
R57 out_buff.n18 out_buff.n0 0.582399
R58 out_buff.n15 out_buff.n11 0.582399
R59 out_buff.n14 out_buff.n12 0.582399
R60 out_buff.n16 out_buff.n10 0.579923
R61 out_buff.n17 out_buff.n16 0.333833
R62 out_buff.n19 out_buff.n18 0.250559
R63 out_buff out_buff.n30 0.05675
R64 gnd.n267 gnd.n264 10830.8
R65 gnd.n137 gnd.n136 6386.79
R66 gnd.n61 gnd.t18 2974.74
R67 gnd.n140 gnd.n137 1867.45
R68 gnd.n137 gnd.t129 1351.39
R69 gnd.n45 gnd.n44 1273.6
R70 gnd.n58 gnd.n57 1260.8
R71 gnd.n54 gnd.n41 1088.88
R72 gnd.n31 gnd.n30 942.902
R73 gnd gnd.n61 644.029
R74 gnd.n206 gnd.n205 585
R75 gnd.n260 gnd.n259 585
R76 gnd.n262 gnd.n261 585
R77 gnd.n165 gnd.n164 585
R78 gnd.n148 gnd.n147 533.923
R79 gnd.t8 gnd.t80 523.77
R80 gnd.n148 gnd.n3 505.849
R81 gnd.n170 gnd.t85 398.539
R82 gnd.n269 gnd.t83 394.255
R83 gnd.t11 gnd.n207 355.685
R84 gnd.t129 gnd.t6 278.673
R85 gnd.t6 gnd.t82 278.673
R86 gnd.t82 gnd.t26 278.673
R87 gnd.t26 gnd.t7 278.673
R88 gnd.t87 gnd.t113 278.673
R89 gnd.t80 gnd.t87 278.673
R90 gnd.t17 gnd.t8 278.673
R91 gnd.t27 gnd.t17 278.673
R92 gnd.t131 gnd.t27 278.673
R93 gnd.t78 gnd.t131 278.673
R94 gnd.t95 gnd.t78 278.673
R95 gnd.t18 gnd.t30 278.673
R96 gnd.t30 gnd.n4 271.957
R97 gnd.n62 gnd.t22 266.197
R98 gnd.n236 gnd.t13 265.693
R99 gnd.n158 gnd.n148 257.24
R100 gnd.t28 gnd.t2 247.738
R101 gnd.n79 gnd.t29 215.036
R102 gnd.t151 gnd.n169 205.698
R103 gnd.t123 gnd.t127 182.645
R104 gnd.t127 gnd.t81 182.645
R105 gnd.n61 gnd.n60 182.377
R106 gnd.n169 gnd.n168 181.058
R107 gnd.n63 gnd.n62 180.341
R108 gnd.n238 gnd.n235 163.766
R109 gnd.t79 gnd.t32 161.273
R110 gnd.n271 gnd.n260 156.236
R111 gnd.n89 gnd.t128 154.317
R112 gnd.n217 gnd.n216 153.976
R113 gnd.n214 gnd.t0 152.131
R114 gnd.t147 gnd.n268 152.131
R115 gnd.n215 gnd.n210 150.648
R116 gnd.n69 gnd.n65 149.835
R117 gnd.t130 gnd.t58 148.88
R118 gnd.t102 gnd.t56 148.88
R119 gnd.t36 gnd.t66 148.88
R120 gnd.t15 gnd.t37 148.88
R121 gnd.t105 gnd.t76 148.88
R122 gnd.t97 gnd.t74 148.88
R123 gnd.t119 gnd.t41 148.88
R124 gnd.t110 gnd.t54 148.88
R125 gnd.t99 gnd.t68 148.88
R126 gnd.t19 gnd.t43 148.88
R127 gnd.t16 gnd.t39 148.88
R128 gnd.t98 gnd.t52 148.88
R129 gnd.t104 gnd.t48 148.88
R130 gnd.t135 gnd.t64 148.88
R131 gnd.n217 gnd.n206 148.707
R132 gnd.t121 gnd.t125 144.756
R133 gnd.n236 gnd.t20 141.417
R134 gnd.t106 gnd.n38 134.613
R135 gnd.n268 gnd.n267 131.775
R136 gnd.n91 gnd.n90 128.757
R137 gnd.t90 gnd.t136 128.24
R138 gnd.n87 gnd.n86 116.754
R139 gnd.n118 gnd.n77 107.24
R140 gnd.n105 gnd.n83 107.24
R141 gnd.t5 gnd.t31 105.895
R142 gnd.n55 gnd.t50 104.216
R143 gnd.t62 gnd.n49 102.975
R144 gnd.t111 gnd.t135 101.734
R145 gnd.t9 gnd.t25 101.734
R146 gnd.n86 gnd.t122 100.001
R147 gnd.n70 gnd.n69 98.6358
R148 gnd.t31 gnd.t90 96.1807
R149 gnd.n208 gnd.t11 94.2786
R150 gnd.t22 gnd.t123 94.2376
R151 gnd.t125 gnd.t5 93.2661
R152 gnd.t32 gnd.t4 93.2661
R153 gnd.t4 gnd.t28 92.2946
R154 gnd.n52 gnd.t46 89.328
R155 gnd.n35 gnd.n34 88.7077
R156 gnd.t81 gnd.t121 88.4085
R157 gnd.n57 gnd.n54 88.0946
R158 gnd.n42 gnd.t60 86.2264
R159 gnd.n39 gnd.t132 81.884
R160 gnd.t2 gnd.t34 81.6079
R161 gnd.t83 gnd.n263 77.1371
R162 gnd.n42 gnd.t45 73.8198
R163 gnd.n83 gnd.t137 72.8576
R164 gnd.n86 gnd.t126 70.0005
R165 gnd.t136 gnd.t79 69.9497
R166 gnd.n172 gnd.n165 65.8829
R167 gnd.t34 gnd 63.1491
R168 gnd.n83 gnd.t91 60.5809
R169 gnd.n41 gnd.n37 60.3613
R170 gnd.n52 gnd.t101 59.5522
R171 gnd.t25 gnd.t111 58.3115
R172 gnd.t103 gnd.t9 58.3115
R173 gnd.n90 gnd.t124 57.1434
R174 gnd.n34 gnd.n31 49.6269
R175 gnd.n271 gnd.n262 48.5652
R176 gnd.n49 gnd.t138 45.9049
R177 gnd.n77 gnd.t3 38.5719
R178 gnd.n77 gnd.t35 38.5719
R179 gnd.n252 gnd.t146 37.3602
R180 gnd.n255 gnd.t169 37.3602
R181 gnd.n258 gnd.t154 37.3602
R182 gnd.n177 gnd.t163 37.3602
R183 gnd.n180 gnd.t157 37.3602
R184 gnd.n183 gnd.t166 37.3602
R185 gnd.n107 gnd.n106 34.6358
R186 gnd.n107 gnd.n81 34.6358
R187 gnd.n111 gnd.n81 34.6358
R188 gnd.n112 gnd.n111 34.6358
R189 gnd.n113 gnd.n112 34.6358
R190 gnd.n99 gnd.n98 34.6358
R191 gnd.n100 gnd.n99 34.6358
R192 gnd.n100 gnd.n84 34.6358
R193 gnd.n104 gnd.n84 34.6358
R194 gnd.n94 gnd.n93 34.6358
R195 gnd.n95 gnd.n94 34.6358
R196 gnd.n117 gnd.n79 29.7417
R197 gnd.n93 gnd.n89 27.8593
R198 gnd.n214 gnd.n211 27.8554
R199 gnd.n90 gnd.t23 25.4291
R200 gnd.n158 gnd.t107 25.1825
R201 gnd.n155 gnd.n152 24.9897
R202 gnd.n119 gnd.n118 24.4919
R203 gnd.t24 gnd.n140 23.5887
R204 gnd.n147 gnd.t24 23.5887
R205 gnd.n118 gnd.n117 22.9652
R206 gnd.n39 gnd.t103 19.8511
R207 gnd.n174 gnd.t150 18.6812
R208 gnd.n249 gnd.t160 18.6809
R209 gnd.n95 gnd.n87 17.6946
R210 gnd.n232 gnd.t144 17.4089
R211 gnd.n202 gnd.t116 17.4089
R212 gnd.n243 gnd.t115 17.4084
R213 gnd.n241 gnd.t84 17.4084
R214 gnd.n240 gnd.t140 17.4084
R215 gnd.n243 gnd.t88 17.4084
R216 gnd.n241 gnd.t114 17.4084
R217 gnd.n240 gnd.t133 17.4084
R218 gnd.n232 gnd.t143 17.4079
R219 gnd.n202 gnd.t96 17.4079
R220 gnd.n245 gnd.t21 17.4074
R221 gnd.n245 gnd.t139 17.4074
R222 gnd.n219 gnd.t117 17.4069
R223 gnd.n219 gnd.t1 17.4055
R224 gnd.n248 gnd.t162 17.405
R225 gnd.n248 gnd.t161 17.405
R226 gnd.n251 gnd.t149 17.405
R227 gnd.n251 gnd.t148 17.405
R228 gnd.n254 gnd.t171 17.405
R229 gnd.n254 gnd.t170 17.405
R230 gnd.n257 gnd.t156 17.405
R231 gnd.n257 gnd.t155 17.405
R232 gnd.n173 gnd.t153 17.405
R233 gnd.n173 gnd.t152 17.405
R234 gnd.n176 gnd.t165 17.405
R235 gnd.n176 gnd.t164 17.405
R236 gnd.n179 gnd.t159 17.405
R237 gnd.n179 gnd.t158 17.405
R238 gnd.n182 gnd.t168 17.405
R239 gnd.n182 gnd.t167 17.405
R240 gnd.n73 gnd.t94 17.405
R241 gnd.n221 gnd.t142 17.4034
R242 gnd.n220 gnd.t14 17.4034
R243 gnd.n227 gnd.t109 17.4034
R244 gnd.n226 gnd.t134 17.4034
R245 gnd.n197 gnd.t86 17.4034
R246 gnd.n196 gnd.t12 17.4034
R247 gnd.n191 gnd.t145 17.4034
R248 gnd.n190 gnd.t141 17.4034
R249 gnd.n186 gnd.t89 17.4034
R250 gnd.n185 gnd.t33 17.4034
R251 gnd.n24 gnd.t112 17.4005
R252 gnd.n24 gnd.t10 17.4005
R253 gnd.n22 gnd.t49 17.4005
R254 gnd.n22 gnd.t65 17.4005
R255 gnd.n20 gnd.t40 17.4005
R256 gnd.n20 gnd.t53 17.4005
R257 gnd.n18 gnd.t69 17.4005
R258 gnd.n18 gnd.t44 17.4005
R259 gnd.n16 gnd.t73 17.4005
R260 gnd.n16 gnd.t71 17.4005
R261 gnd.n14 gnd.t47 17.4005
R262 gnd.n14 gnd.t63 17.4005
R263 gnd.n12 gnd.t55 17.4005
R264 gnd.n12 gnd.t51 17.4005
R265 gnd.n10 gnd.t75 17.4005
R266 gnd.n10 gnd.t42 17.4005
R267 gnd.n8 gnd.t38 17.4005
R268 gnd.n8 gnd.t77 17.4005
R269 gnd.n6 gnd.t57 17.4005
R270 gnd.n6 gnd.t67 17.4005
R271 gnd.n5 gnd.t61 17.4005
R272 gnd.n5 gnd.t59 17.4005
R273 gnd.n113 gnd.n79 14.6829
R274 gnd.n38 gnd.t70 14.2681
R275 gnd.n269 gnd.t147 12.8566
R276 gnd.t56 gnd.t130 11.1664
R277 gnd.t66 gnd.t102 11.1664
R278 gnd.t37 gnd.t36 11.1664
R279 gnd.t76 gnd.t15 11.1664
R280 gnd.t74 gnd.t105 11.1664
R281 gnd.t41 gnd.t97 11.1664
R282 gnd.t54 gnd.t119 11.1664
R283 gnd.t50 gnd.t110 11.1664
R284 gnd.t46 gnd.t100 11.1664
R285 gnd.t101 gnd.t62 11.1664
R286 gnd.t138 gnd.t72 11.1664
R287 gnd.t70 gnd.t120 11.1664
R288 gnd.t68 gnd.t106 11.1664
R289 gnd.t43 gnd.t99 11.1664
R290 gnd.t39 gnd.t19 11.1664
R291 gnd.t52 gnd.t16 11.1664
R292 gnd.t48 gnd.t98 11.1664
R293 gnd.t64 gnd.t104 11.1664
R294 gnd.n91 gnd.n89 10.9075
R295 gnd.n73 gnd.n72 9.33321
R296 gnd.n172 gnd.n171 9.3005
R297 gnd.n171 gnd.n170 9.3005
R298 gnd.n217 gnd.n209 9.3005
R299 gnd.n209 gnd.n208 9.3005
R300 gnd.n238 gnd.n237 9.3005
R301 gnd.n237 gnd.n236 9.3005
R302 gnd.n271 gnd.n270 9.3005
R303 gnd.n270 gnd.n269 9.3005
R304 gnd.n162 gnd.t108 8.70236
R305 gnd.n170 gnd.t151 8.57123
R306 gnd.n106 gnd.n105 7.90638
R307 gnd.n4 gnd.t95 6.71549
R308 gnd.n35 gnd.t118 4.96314
R309 gnd.n115 gnd.n79 4.6505
R310 gnd.n93 gnd.n92 4.6505
R311 gnd.n94 gnd.n88 4.6505
R312 gnd.n96 gnd.n95 4.6505
R313 gnd.n98 gnd.n97 4.6505
R314 gnd.n99 gnd.n85 4.6505
R315 gnd.n101 gnd.n100 4.6505
R316 gnd.n102 gnd.n84 4.6505
R317 gnd.n104 gnd.n103 4.6505
R318 gnd.n106 gnd.n82 4.6505
R319 gnd.n108 gnd.n107 4.6505
R320 gnd.n109 gnd.n81 4.6505
R321 gnd.n111 gnd.n110 4.6505
R322 gnd.n112 gnd.n80 4.6505
R323 gnd.n114 gnd.n113 4.6505
R324 gnd.n117 gnd.n116 4.6505
R325 gnd.n118 gnd.n78 4.6505
R326 gnd.n75 gnd.n74 4.5005
R327 gnd.n76 gnd.n74 4.5005
R328 gnd gnd.n122 3.79922
R329 gnd.n123 gnd.n0 3.24248
R330 gnd.n26 gnd.n0 3.01925
R331 gnd.n126 gnd.n124 2.6505
R332 gnd.n98 gnd.n87 2.63579
R333 gnd gnd.n162 2.5773
R334 gnd.n120 gnd.n74 2.25328
R335 gnd.n105 gnd.n104 1.88285
R336 gnd.n163 gnd 1.8224
R337 gnd.n7 gnd.n5 1.66573
R338 gnd.n124 gnd.t92 1.47915
R339 gnd.n25 gnd.n23 1.3755
R340 gnd.n163 gnd.n0 1.30732
R341 gnd.n124 gnd.n123 1.22706
R342 gnd.n9 gnd.n7 1.08383
R343 gnd.n13 gnd.n11 1.08383
R344 gnd.n15 gnd.n13 1.08383
R345 gnd.n17 gnd.n15 1.08383
R346 gnd.n21 gnd.n19 1.08383
R347 gnd.n23 gnd.n21 1.08383
R348 gnd.n11 gnd.n9 1.04217
R349 gnd.n19 gnd.n17 1.04217
R350 gnd.n23 gnd.n22 0.582399
R351 gnd.n21 gnd.n20 0.582399
R352 gnd.n19 gnd.n18 0.582399
R353 gnd.n17 gnd.n16 0.582399
R354 gnd.n15 gnd.n14 0.582399
R355 gnd.n13 gnd.n12 0.582399
R356 gnd.n11 gnd.n10 0.582399
R357 gnd.n7 gnd.n6 0.582399
R358 gnd.n9 gnd.n8 0.579923
R359 gnd.n25 gnd.n24 0.57713
R360 gnd.n130 gnd.n71 0.54125
R361 gnd.n71 gnd.n70 0.541165
R362 gnd.n225 gnd.n219 0.447415
R363 gnd.n231 gnd.n225 0.438
R364 gnd.n233 gnd.n231 0.438
R365 gnd.n275 gnd.n274 0.401236
R366 gnd.n27 gnd.n25 0.392443
R367 gnd.n195 gnd.n189 0.375501
R368 gnd.n234 gnd.n233 0.375501
R369 gnd.n201 gnd.n195 0.3755
R370 gnd.n203 gnd.n201 0.3755
R371 gnd.n242 gnd.n240 0.373217
R372 gnd.n244 gnd.n242 0.371401
R373 gnd.n246 gnd.n244 0.369555
R374 gnd.n159 gnd.n2 0.366293
R375 gnd.n150 gnd.n149 0.365897
R376 gnd.n158 gnd.n150 0.365897
R377 gnd.n2 gnd.n1 0.365897
R378 gnd.n135 gnd.n134 0.347558
R379 gnd.n134 gnd.n133 0.347269
R380 gnd.n247 gnd.n246 0.338503
R381 gnd.n204 gnd.n203 0.330858
R382 gnd.n204 gnd.n184 0.290469
R383 gnd.n37 gnd.n36 0.288252
R384 gnd.n36 gnd.n35 0.288252
R385 gnd.n234 gnd.n218 0.281539
R386 gnd.n27 gnd.n26 0.274914
R387 gnd.n239 gnd.n234 0.245825
R388 gnd.n273 gnd.n247 0.244548
R389 gnd.n275 gnd.n163 0.230614
R390 gnd.n247 gnd.n239 0.180349
R391 gnd.n218 gnd.n204 0.156539
R392 gnd.n92 gnd.n91 0.144332
R393 gnd.n142 gnd.n141 0.1305
R394 gnd.t24 gnd.n142 0.1305
R395 gnd.n144 gnd.n143 0.1305
R396 gnd.t24 gnd.n144 0.1305
R397 gnd.n92 gnd.n88 0.120292
R398 gnd.n96 gnd.n88 0.120292
R399 gnd.n97 gnd.n96 0.120292
R400 gnd.n97 gnd.n85 0.120292
R401 gnd.n101 gnd.n85 0.120292
R402 gnd.n102 gnd.n101 0.120292
R403 gnd.n103 gnd.n102 0.120292
R404 gnd.n103 gnd.n82 0.120292
R405 gnd.n108 gnd.n82 0.120292
R406 gnd.n109 gnd.n108 0.120292
R407 gnd.n110 gnd.n109 0.120292
R408 gnd.n110 gnd.n80 0.120292
R409 gnd.n114 gnd.n80 0.120292
R410 gnd.n115 gnd.n114 0.120292
R411 gnd.n116 gnd.n115 0.120292
R412 gnd.n116 gnd.n78 0.120292
R413 gnd.n154 gnd.n153 0.10956
R414 gnd.n157 gnd.n156 0.10956
R415 gnd.t107 gnd.n157 0.10956
R416 gnd.n67 gnd.n66 0.10956
R417 gnd.t93 gnd.n67 0.10956
R418 gnd.n68 gnd.t93 0.10956
R419 gnd.n69 gnd.n68 0.10956
R420 gnd.n155 gnd.n154 0.109112
R421 gnd.n135 gnd.n132 0.0849523
R422 gnd.n132 gnd.n131 0.0845034
R423 gnd.n276 gnd.n275 0.0772045
R424 gnd.n276 gnd 0.0755
R425 gnd.n78 gnd.n75 0.0734167
R426 gnd.n250 gnd.n249 0.073412
R427 gnd.n175 gnd.n174 0.0734113
R428 gnd.n26 gnd 0.06925
R429 gnd.n176 gnd.n175 0.0610469
R430 gnd.n177 gnd.n176 0.0610469
R431 gnd.n179 gnd.n178 0.0610469
R432 gnd.n180 gnd.n179 0.0610469
R433 gnd.n182 gnd.n181 0.0610469
R434 gnd.n183 gnd.n182 0.0610469
R435 gnd.n251 gnd.n250 0.0610469
R436 gnd.n252 gnd.n251 0.0610469
R437 gnd.n254 gnd.n253 0.0610469
R438 gnd.n255 gnd.n254 0.0610469
R439 gnd.n257 gnd.n256 0.0610469
R440 gnd.n258 gnd.n257 0.0610469
R441 gnd.n272 gnd.n258 0.0573558
R442 gnd.n184 gnd.n183 0.0573547
R443 gnd.n273 gnd.n272 0.0464211
R444 gnd.n178 gnd.n177 0.0426875
R445 gnd.n181 gnd.n180 0.0426875
R446 gnd.n253 gnd.n252 0.0426875
R447 gnd.n256 gnd.n255 0.0426875
R448 gnd.n65 gnd.n64 0.0425017
R449 gnd.n64 gnd.n63 0.0425017
R450 gnd.n29 gnd.n28 0.0425017
R451 gnd.n31 gnd.n29 0.0425017
R452 gnd.n44 gnd.n43 0.0425017
R453 gnd.n43 gnd.n42 0.0425017
R454 gnd.n33 gnd.n32 0.0425017
R455 gnd.n34 gnd.n33 0.0425017
R456 gnd.n59 gnd.n58 0.0425017
R457 gnd.n60 gnd.n59 0.0425017
R458 gnd.n274 gnd 0.0395625
R459 gnd gnd.n276 0.0345909
R460 gnd.n76 gnd 0.0330521
R461 gnd.n123 gnd 0.03175
R462 gnd.n174 gnd.n173 0.031274
R463 gnd.n249 gnd.n248 0.0312734
R464 gnd.n121 gnd.n75 0.0265417
R465 gnd.n152 gnd.n151 0.0264102
R466 gnd.n119 gnd 0.0226354
R467 gnd.n233 gnd.n232 0.0153409
R468 gnd.n230 gnd.n228 0.0129048
R469 gnd.n121 gnd.n120 0.0114272
R470 gnd.n224 gnd.n222 0.0114167
R471 gnd.n120 gnd.n119 0.0113582
R472 gnd.n122 gnd.n74 0.0110001
R473 gnd.n216 gnd.n215 0.0092427
R474 gnd.n215 gnd.n214 0.0092427
R475 gnd.n266 gnd.n265 0.00883856
R476 gnd.n267 gnd.n266 0.00883856
R477 gnd.n167 gnd.n166 0.00883856
R478 gnd.n168 gnd.n167 0.00883856
R479 gnd.n127 gnd.n73 0.00867757
R480 gnd.n203 gnd.n202 0.00792873
R481 gnd.n146 gnd.n145 0.00762598
R482 gnd.n147 gnd.n146 0.00762598
R483 gnd.n139 gnd.n138 0.00762598
R484 gnd.n140 gnd.n139 0.00762598
R485 gnd.n127 gnd.n126 0.00634112
R486 gnd gnd.n76 0.00570833
R487 gnd.n200 gnd.n198 0.00546432
R488 gnd.n187 gnd.n185 0.00502806
R489 gnd.n192 gnd.n190 0.00502806
R490 gnd.n198 gnd.n196 0.00502805
R491 gnd.n222 gnd.n220 0.00502803
R492 gnd.n228 gnd.n226 0.00502803
R493 gnd.n57 gnd.n56 0.00498892
R494 gnd.n56 gnd.n55 0.00498892
R495 gnd.n213 gnd.n212 0.00487141
R496 gnd.n214 gnd.n213 0.00487141
R497 gnd.n54 gnd.n53 0.00466542
R498 gnd.n53 gnd.n52 0.00466542
R499 gnd.n130 gnd.n129 0.00441022
R500 gnd.n187 gnd.n186 0.00402807
R501 gnd.n192 gnd.n191 0.00402806
R502 gnd.n198 gnd.n197 0.00402806
R503 gnd.n222 gnd.n221 0.00402804
R504 gnd.n228 gnd.n227 0.00402803
R505 gnd.n194 gnd.n192 0.00397623
R506 gnd.n129 gnd.n128 0.00391284
R507 gnd.n128 gnd.n127 0.00391159
R508 gnd.n46 gnd.n45 0.00271942
R509 gnd.n49 gnd.n46 0.00271942
R510 gnd.n48 gnd.n47 0.00271942
R511 gnd.n49 gnd.n48 0.00271942
R512 gnd.n51 gnd.n50 0.00258271
R513 gnd.n52 gnd.n51 0.00258271
R514 gnd.n189 gnd.n187 0.00248813
R515 gnd.n274 gnd.n273 0.00245312
R516 gnd.n160 gnd.n159 0.00236777
R517 gnd.t107 gnd.n155 0.00194448
R518 gnd.n41 gnd.n40 0.00190526
R519 gnd.n40 gnd.n39 0.00190526
R520 gnd.n161 gnd.n160 0.00186816
R521 gnd.n272 gnd.n271 0.00152216
R522 gnd.n184 gnd.n172 0.00152195
R523 gnd.n230 gnd.n229 0.00138337
R524 gnd.n224 gnd.n223 0.00138109
R525 gnd.n200 gnd.n199 0.00134613
R526 gnd.n194 gnd.n193 0.00134049
R527 gnd.n189 gnd.n188 0.001335
R528 gnd.n162 gnd.n161 0.00124275
R529 gnd.n244 gnd.n243 0.00121065
R530 gnd.n242 gnd.n241 0.001204
R531 gnd.n136 gnd.n135 0.00104118
R532 gnd.n122 gnd.n121 0.00100955
R533 gnd.n136 gnd.n130 0.00100261
R534 gnd.n246 gnd.n245 0.00100079
R535 gnd.n159 gnd.n158 0.00100039
R536 gnd.n218 gnd.n217 0.000522345
R537 gnd.n239 gnd.n238 0.000522345
R538 gnd.n126 gnd.n125 0.00051897
R539 gnd.n41 gnd.n27 0.000503131
R540 gnd.n231 gnd.n230 0.000501021
R541 gnd.n225 gnd.n224 0.000501021
R542 gnd.n195 gnd.n194 0.000500672
R543 gnd.n201 gnd.n200 0.000500672
R544 buffer_0.a.n6 buffer_0.a.t26 40.2461
R545 buffer_0.a.n2 buffer_0.a.t21 40.2461
R546 buffer_0.a.n10 buffer_0.a.t5 39.5292
R547 buffer_0.a.n9 buffer_0.a.t20 39.5292
R548 buffer_0.a.n8 buffer_0.a.t17 39.5292
R549 buffer_0.a.n7 buffer_0.a.t25 39.5292
R550 buffer_0.a.n6 buffer_0.a.t18 39.5292
R551 buffer_0.a.n5 buffer_0.a.t19 39.5292
R552 buffer_0.a.n4 buffer_0.a.t24 39.5292
R553 buffer_0.a.n3 buffer_0.a.t23 39.5292
R554 buffer_0.a.n2 buffer_0.a.t22 39.5292
R555 buffer_0.a.n12 buffer_0.a.t6 28.576
R556 buffer_0.a.n1 buffer_0.a.t2 25.2845
R557 buffer_0.a.n0 buffer_0.a.t0 24.699
R558 buffer_0.a.n1 buffer_0.a.t4 17.4081
R559 buffer_0.a.n1 buffer_0.a.t9 17.4005
R560 buffer_0.a.n1 buffer_0.a.t3 17.4005
R561 buffer_0.a.n17 buffer_0.a.t16 17.4005
R562 buffer_0.a.n17 buffer_0.a.t14 17.4005
R563 buffer_0.a.n15 buffer_0.a.t11 17.4005
R564 buffer_0.a.n15 buffer_0.a.t10 17.4005
R565 buffer_0.a.n13 buffer_0.a.t15 17.4005
R566 buffer_0.a.n13 buffer_0.a.t12 17.4005
R567 buffer_0.a.n0 buffer_0.a.t1 17.4005
R568 buffer_0.a.n0 buffer_0.a.t13 17.4005
R569 buffer_0.a.n19 buffer_0.a.t7 17.4005
R570 buffer_0.a.n19 buffer_0.a.t8 17.4005
R571 buffer_0.a.n14 buffer_0.a.n0 2.76905
R572 buffer_0.a.n20 buffer_0.a.n1 2.69153
R573 buffer_0.a.n16 buffer_0.a.n14 2.16717
R574 buffer_0.a.n18 buffer_0.a.n16 2.1255
R575 buffer_0.a.n21 buffer_0.a.n20 1.2505
R576 buffer_0.a.n10 buffer_0.a.n9 1.06739
R577 buffer_0.a.n21 buffer_0.a.n18 0.917167
R578 buffer_0.a buffer_0.a.n12 0.862147
R579 buffer_0.a.n11 buffer_0.a.n5 0.749569
R580 buffer_0.a.n7 buffer_0.a.n6 0.717388
R581 buffer_0.a.n8 buffer_0.a.n7 0.717388
R582 buffer_0.a.n9 buffer_0.a.n8 0.717388
R583 buffer_0.a.n3 buffer_0.a.n2 0.717388
R584 buffer_0.a.n4 buffer_0.a.n3 0.717388
R585 buffer_0.a.n5 buffer_0.a.n4 0.717388
R586 buffer_0.a.n20 buffer_0.a.n19 0.526026
R587 buffer_0.a.n16 buffer_0.a.n15 0.52595
R588 buffer_0.a buffer_0.a.n21 0.521392
R589 buffer_0.a.n18 buffer_0.a.n17 0.516495
R590 buffer_0.a.n14 buffer_0.a.n13 0.516495
R591 buffer_0.a.n11 buffer_0.a.n10 0.349569
R592 buffer_0.a.n12 buffer_0.a.n11 0.271856
R593 vd.n62 vd.n59 2142.35
R594 vd.n31 vd.n28 1304.47
R595 vd.n66 vd.n60 1164.71
R596 vd.n68 vd.n56 1164.71
R597 vd.n44 vd.n36 1070.68
R598 vd.n68 vd.n57 977.648
R599 vd.n66 vd.n59 952.942
R600 vd.t63 vd.t73 537.318
R601 vd.t73 vd.t75 526.24
R602 vd.t15 vd.t17 526.24
R603 vd.t13 vd.t15 512.391
R604 vd.t54 vd.t77 357.289
R605 vd.t77 vd.t65 357.289
R606 vd.t65 vd.t61 357.289
R607 vd.t75 vd.t57 357.289
R608 vd.t59 vd.t63 357.289
R609 vd.t69 vd.t59 357.289
R610 vd.t67 vd.t69 357.289
R611 vd.t11 vd.t9 357.289
R612 vd.t9 vd.t7 357.289
R613 vd.t7 vd.t5 357.289
R614 vd.t21 vd.t13 357.289
R615 vd.t3 vd.t21 357.289
R616 vd.t19 vd.t3 357.289
R617 vd.n27 vd.t54 354.529
R618 vd.n34 vd.t11 282.507
R619 vd.n34 vd.t71 254.811
R620 vd.n64 vd.n63 228.518
R621 vd.n63 vd.n54 228.518
R622 vd.n43 vd.n40 223.625
R623 vd.n128 vd.n125 206.306
R624 vd.n37 vd.t1 204.957
R625 vd.n96 vd.n95 168.66
R626 vd.t38 vd.n109 156.245
R627 vd.n37 vd.t19 152.333
R628 vd.n67 vd.t32 144.606
R629 vd.n29 vd.t67 144.024
R630 vd.n91 vd.t82 143.697
R631 vd.n113 vd.t30 143.697
R632 vd.n135 vd.n132 142.306
R633 vd.n62 vd.n61 135.465
R634 vd.n36 vd.n31 127.248
R635 vd.n115 vd.n112 126.871
R636 vd.n44 vd.n43 117.835
R637 vd.n88 vd.n87 111.421
R638 vd.n69 vd.n54 104.282
R639 vd.n65 vd.n64 101.647
R640 vd.n41 vd.t46 92.7848
R641 vd.n133 vd.t23 86.6752
R642 vd.n96 vd.n90 85.0829
R643 vd.n126 vd.t42 71.8492
R644 vd.n91 vd.t50 65.0065
R645 vd.n84 vd.t49 63.6934
R646 vd.n98 vd.t41 63.6821
R647 vd.n104 vd.t37 63.6292
R648 vd.n128 vd.n122 63.2476
R649 vd.n133 vd.t79 60.4447
R650 vd.t23 vd.t24 58.1638
R651 vd.t42 vd.t26 58.1638
R652 vd.n120 vd.t27 42.1974
R653 vd.n123 vd.t81 42.1974
R654 vd.n70 vd.n69 31.105
R655 vd.n20 vd.t16 29.2512
R656 vd.n15 vd.t12 29.2303
R657 vd.n10 vd.t64 29.2303
R658 vd.n9 vd.t74 29.2303
R659 vd.n26 vd.t48 28.5795
R660 vd.n3 vd.t78 28.57
R661 vd.n23 vd.t4 28.5655
R662 vd.n23 vd.t20 28.5655
R663 vd.n21 vd.t14 28.5655
R664 vd.n21 vd.t22 28.5655
R665 vd.n18 vd.t6 28.5655
R666 vd.n18 vd.t18 28.5655
R667 vd.n16 vd.t10 28.5655
R668 vd.n16 vd.t8 28.5655
R669 vd.n13 vd.t68 28.5655
R670 vd.n13 vd.t72 28.5655
R671 vd.n11 vd.t60 28.5655
R672 vd.n11 vd.t70 28.5655
R673 vd.n7 vd.t58 28.5655
R674 vd.n7 vd.t76 28.5655
R675 vd.n5 vd.t66 28.5655
R676 vd.n5 vd.t62 28.5655
R677 vd.n25 vd.t2 28.5655
R678 vd.n25 vd.t47 28.5655
R679 vd.n93 vd.t36 28.5119
R680 vd.n65 vd.n48 27.9188
R681 vd.n106 vd.n101 24.5501
R682 vd.n70 vd.n53 22.401
R683 vd.n78 vd.n77 22.4005
R684 vd.n53 vd.n51 22.4005
R685 vd.n110 vd.t38 21.0989
R686 vd.n4 vd.t53 19.8115
R687 vd.n26 vd.t45 19.8115
R688 vd.t27 vd.t29 19.3883
R689 vd.n79 vd.n48 19.201
R690 vd.n79 vd.n78 19.2005
R691 vd.n126 vd.t56 17.1073
R692 vd.n97 vd.t28 14.5056
R693 vd.n83 vd.t25 14.472
R694 vd.n97 vd.t43 14.4415
R695 vd.n99 vd.t44 14.4153
R696 vd.n85 vd.t51 14.4127
R697 vd.n103 vd.t39 14.4041
R698 vd.n83 vd.t52 14.3878
R699 vd.n101 vd.t40 14.2867
R700 vd.n3 vd.t55 14.2847
R701 vd.n102 vd.t31 14.283
R702 vd.n102 vd.t35 14.283
R703 vd.t50 vd.t80 11.4051
R704 vd.n55 vd.n51 10.5605
R705 vd.n77 vd.n50 9.6005
R706 vd.n2 vd.t0 9.5742
R707 vd.n74 vd.t33 9.52337
R708 vd.n106 vd.n105 9.3005
R709 vd.n107 vd.n106 4.5005
R710 vd.n141 vd.n140 3.73002
R711 vd.n113 vd.t34 3.42187
R712 vd vd.n82 2.438
R713 vd.n55 vd.n50 2.2405
R714 vd.n139 vd 2.08242
R715 vd vd.n107 1.83279
R716 vd.n6 vd.n4 1.47391
R717 vd vd.n26 1.0363
R718 vd.n9 vd.n8 1.0005
R719 vd.n20 vd.n19 1.0005
R720 vd.n138 vd.n85 0.862412
R721 vd.n139 vd.n138 0.834744
R722 vd.n8 vd.n6 0.813
R723 vd.n12 vd.n10 0.813
R724 vd.n19 vd.n17 0.813
R725 vd.n14 vd.n12 0.78175
R726 vd.n17 vd.n15 0.78175
R727 vd.n24 vd.n22 0.78175
R728 vd.n103 vd.n102 0.721906
R729 vd.n24 vd.n23 0.665316
R730 vd.n22 vd.n21 0.665316
R731 vd.n19 vd.n18 0.665316
R732 vd.n14 vd.n13 0.665316
R733 vd.n12 vd.n11 0.665316
R734 vd.n8 vd.n7 0.665316
R735 vd.n6 vd.n5 0.665316
R736 vd.n15 vd.n14 0.6255
R737 vd.n17 vd.n16 0.611443
R738 vd.n104 vd.n103 0.608294
R739 vd.n22 vd.n20 0.59425
R740 vd.n117 vd.n99 0.576317
R741 vd.n137 vd.n136 0.5755
R742 vd.n136 vd.n129 0.488
R743 vd.n117 vd.n116 0.463
R744 vd.n99 vd.n98 0.344245
R745 vd.n46 vd.n24 0.302583
R746 vd.n116 vd 0.2755
R747 vd.n129 vd.n117 0.238
R748 vd.n140 vd.n46 0.23013
R749 vd.n10 vd.n9 0.21925
R750 vd.n142 vd.n141 0.2005
R751 vd.n72 vd.n71 0.146341
R752 vd.n72 vd.n47 0.146333
R753 vd.n66 vd.n65 0.130052
R754 vd.n67 vd.n66 0.130052
R755 vd.n84 vd.n83 0.129979
R756 vd.n82 vd.n47 0.1255
R757 vd.n142 vd 0.1255
R758 vd.n101 vd.n100 0.122252
R759 vd.n105 vd.n104 0.116172
R760 vd.n69 vd.n68 0.107375
R761 vd.n68 vd.n67 0.107375
R762 vd.n142 vd.n2 0.0822638
R763 vd.n0 vd.t83 0.0686501
R764 vd.n1 vd.n0 0.06865
R765 vd.n140 vd.n139 0.0648158
R766 vd.n76 vd.n49 0.0456031
R767 vd.n73 vd.n52 0.0456031
R768 vd.n71 vd.n52 0.0456031
R769 vd.n45 vd 0.0421667
R770 vd.n81 vd.n80 0.0391598
R771 vd.n80 vd.n49 0.0391598
R772 vd.n141 vd 0.0372647
R773 vd.n64 vd.n59 0.0349892
R774 vd.n59 vd.t32 0.0349892
R775 vd.n57 vd.n54 0.0349892
R776 vd.n61 vd.n57 0.0333079
R777 vd.n98 vd.n97 0.0321654
R778 vd.n90 vd.n89 0.0307238
R779 vd.n89 vd.n88 0.0302348
R780 vd.n85 vd.n84 0.0267443
R781 vd.n74 vd.n73 0.0217629
R782 vd.n76 vd.n75 0.0198299
R783 vd.n107 vd.n100 0.0176875
R784 vd.n112 vd.n111 0.0175052
R785 vd.n111 vd.n110 0.0175052
R786 vd.n43 vd.n42 0.0168558
R787 vd.n42 vd.n41 0.0168558
R788 vd.n132 vd.n131 0.0150968
R789 vd.n131 vd.n130 0.0150968
R790 vd vd.n142 0.013
R791 vd.n58 vd.n56 0.0125538
R792 vd.n95 vd.n94 0.0122827
R793 vd.n94 vd.n93 0.0122827
R794 vd.n56 vd.n55 0.0120596
R795 vd.n46 vd.n45 0.0109167
R796 vd.n105 vd.n100 0.009875
R797 vd.n40 vd.n39 0.00979742
R798 vd.n28 vd.n27 0.00979742
R799 vd.n125 vd.n124 0.00973799
R800 vd.n124 vd.n123 0.00973799
R801 vd.n2 vd.n1 0.00846782
R802 vd.n138 vd.n137 0.00675
R803 vd.n63 vd.n62 0.00627981
R804 vd.n44 vd.n38 0.0055
R805 vd.n38 vd.n37 0.0055
R806 vd.n75 vd.n74 0.00501031
R807 vd.n4 vd.n3 0.00500317
R808 vd.n26 vd.n25 0.00454578
R809 vd.n135 vd.n134 0.00391284
R810 vd.n134 vd.n133 0.00391284
R811 vd.n128 vd.n127 0.00391284
R812 vd.n127 vd.n126 0.00391284
R813 vd.n115 vd.n114 0.00391284
R814 vd.n114 vd.n113 0.00391284
R815 vd.n96 vd.n92 0.00391284
R816 vd.n92 vd.n91 0.00391284
R817 vd.n109 vd.n108 0.00347027
R818 vd.n87 vd.n86 0.00347027
R819 vd.n61 vd.t32 0.00318081
R820 vd.n122 vd.n121 0.00275116
R821 vd.n121 vd.n120 0.00275116
R822 vd.n31 vd.n30 0.00186586
R823 vd.n30 vd.n29 0.00186586
R824 vd.n60 vd.n58 0.0018171
R825 vd.n36 vd.n35 0.00173262
R826 vd.n35 vd.n34 0.00173262
R827 vd.n120 vd.n119 0.00162558
R828 vd.n119 vd.n118 0.00162558
R829 vd.n60 vd.n50 0.00131751
R830 vd.n75 vd.n50 0.00131744
R831 vd.n80 vd.n79 0.00119114
R832 vd.n33 vd.n32 0.00111631
R833 vd.n34 vd.n33 0.00111631
R834 vd.n81 vd.n48 0.00101609
R835 vd.n67 vd.n58 0.00100038
R836 vd.n71 vd.n70 0.00100009
R837 vd.n53 vd.n52 0.000659706
R838 vd.n77 vd.n76 0.000659706
R839 vd.n78 vd.n49 0.000543686
R840 vd.n73 vd.n51 0.000543686
R841 vd.n136 vd.n135 0.000532663
R842 vd.n129 vd.n128 0.000532663
R843 vd.n116 vd.n115 0.000532663
R844 vd.n137 vd.n96 0.000532663
R845 vd.n45 vd.n44 0.000511142
R846 vd.n82 vd.n81 0.000507883
R847 vd.n49 vd.n47 0.000507883
R848 vd.n73 vd.n72 0.000507883
R849 vd.n0 vd.t85 0.000500086
R850 vd.n1 vd.t84 0.000500086
R851 sensor_0.b.t10 sensor_0.b.t2 74.8549
R852 sensor_0.b.t8 sensor_0.b.t10 74.8549
R853 sensor_0.b.t16 sensor_0.b.t8 74.8549
R854 sensor_0.b.t12 sensor_0.b.t4 74.8549
R855 sensor_0.b.t6 sensor_0.b.t12 74.8549
R856 sensor_0.b.t14 sensor_0.b.t6 74.8549
R857 sensor_0.b.t24 sensor_0.b.t32 74.8549
R858 sensor_0.b.t31 sensor_0.b.t24 74.8549
R859 sensor_0.b.t23 sensor_0.b.t31 74.8549
R860 sensor_0.b.t34 sensor_0.b.t26 74.8549
R861 sensor_0.b.t21 sensor_0.b.t34 74.8549
R862 sensor_0.b.t29 sensor_0.b.t21 74.8549
R863 sensor_0.b.t27 sensor_0.b.t20 74.8549
R864 sensor_0.b.t28 sensor_0.b.t27 74.8549
R865 sensor_0.b.t35 sensor_0.b.t28 74.8549
R866 sensor_0.b.t22 sensor_0.b.t30 74.8549
R867 sensor_0.b.t33 sensor_0.b.t22 74.8549
R868 sensor_0.b.t25 sensor_0.b.t33 74.8549
R869 sensor_0.b.n7 sensor_0.b.t25 38.3763
R870 sensor_0.b.n11 sensor_0.b.t16 37.3627
R871 sensor_0.b.n10 sensor_0.b.t14 37.3602
R872 sensor_0.b.n9 sensor_0.b.t23 37.3602
R873 sensor_0.b.n8 sensor_0.b.t29 37.3602
R874 sensor_0.b.n7 sensor_0.b.t35 37.3602
R875 sensor_0.b.n12 sensor_0.b.t3 18.2715
R876 sensor_0.b.n3 sensor_0.b.t5 18.1717
R877 sensor_0.b.n14 sensor_0.b.t17 17.427
R878 sensor_0.b.n13 sensor_0.b.t9 17.4116
R879 sensor_0.b.n3 sensor_0.b.t13 17.4101
R880 sensor_0.b.n12 sensor_0.b.t11 17.4101
R881 sensor_0.b.n4 sensor_0.b.t7 17.4058
R882 sensor_0.b.n5 sensor_0.b.t15 17.4056
R883 sensor_0.b.n0 sensor_0.b.t19 14.283
R884 sensor_0.b.n0 sensor_0.b.t1 14.283
R885 sensor_0.b.n1 sensor_0.b.t0 14.283
R886 sensor_0.b.n1 sensor_0.b.t18 14.283
R887 sensor_0.b.n6 sensor_0.b.n5 3.22928
R888 sensor_0.b.n6 sensor_0.b.n2 2.2255
R889 sensor_0.b.n11 sensor_0.b.n10 1.01759
R890 sensor_0.b.n8 sensor_0.b.n7 1.01657
R891 sensor_0.b.n9 sensor_0.b.n8 1.01657
R892 sensor_0.b.n10 sensor_0.b.n9 1.01657
R893 sensor_0.b.n13 sensor_0.b.n12 0.865287
R894 sensor_0.b sensor_0.b.n15 0.851048
R895 sensor_0.b.n14 sensor_0.b.n13 0.777059
R896 sensor_0.b.n5 sensor_0.b.n4 0.718555
R897 sensor_0.b.n4 sensor_0.b.n3 0.710921
R898 sensor_0.b.n2 sensor_0.b.n0 0.49917
R899 sensor_0.b sensor_0.b.n6 0.341125
R900 sensor_0.b.n15 sensor_0.b.n14 0.325292
R901 sensor_0.b.n15 sensor_0.b.n11 0.202053
R902 sensor_0.b.n2 sensor_0.b.n1 0.17167
R903 sensor_0.a.n2 sensor_0.a.t15 64.1667
R904 sensor_0.a.n0 sensor_0.a.t0 63.6292
R905 sensor_0.a.n4 sensor_0.a.t13 63.6292
R906 sensor_0.a.n3 sensor_0.a.t12 63.6292
R907 sensor_0.a.n2 sensor_0.a.t14 63.6292
R908 sensor_0.a.n1 sensor_0.a.t2 63.6275
R909 sensor_0.a.n8 sensor_0.a.t6 18.2715
R910 sensor_0.a.n5 sensor_0.a.t11 18.2714
R911 sensor_0.a.n10 sensor_0.a.t9 17.4132
R912 sensor_0.a.n7 sensor_0.a.t4 17.4132
R913 sensor_0.a.n6 sensor_0.a.t7 17.4116
R914 sensor_0.a.n8 sensor_0.a.t10 17.4101
R915 sensor_0.a.n5 sensor_0.a.t8 17.4101
R916 sensor_0.a.n9 sensor_0.a.t5 17.4057
R917 sensor_0.a.n1 sensor_0.a.t3 14.5343
R918 sensor_0.a.n0 sensor_0.a.t1 14.2976
R919 sensor_0.a sensor_0.a.n11 1.63801
R920 sensor_0.a.n11 sensor_0.a.n7 1.541
R921 sensor_0.a.n11 sensor_0.a.n10 1.541
R922 sensor_0.a.n10 sensor_0.a.n9 0.873387
R923 sensor_0.a.n6 sensor_0.a.n5 0.865287
R924 sensor_0.a.n7 sensor_0.a.n6 0.864262
R925 sensor_0.a.n9 sensor_0.a.n8 0.848309
R926 sensor_0.a.n3 sensor_0.a.n2 0.538
R927 sensor_0.a.n4 sensor_0.a.n3 0.538
R928 sensor_0.a.n0 sensor_0.a.n4 0.488
R929 sensor_0.a.n1 sensor_0.a.n0 0.29354
R930 sensor_0.a sensor_0.a.n1 0.28675
R931 vpwr.t1 vpwr.t12 790.188
R932 vpwr.t28 vpwr.t24 648.131
R933 vpwr.t8 vpwr.t20 583.023
R934 vpwr.n77 vpwr 548.548
R935 vpwr.n56 vpwr.t21 514.011
R936 vpwr.t18 vpwr.t28 485.358
R937 vpwr.t0 vpwr.t16 414.33
R938 vpwr.n14 vpwr.t7 413.315
R939 vpwr.n32 vpwr.t13 375.277
R940 vpwr.n7 vpwr.t4 344.005
R941 vpwr.t26 vpwr.t5 319.627
R942 vpwr.n50 vpwr.n39 311.957
R943 vpwr.n72 vpwr.n31 311.894
R944 vpwr.n59 vpwr.n58 309.18
R945 vpwr.t20 vpwr.t3 292.991
R946 vpwr.t14 vpwr.t0 292.991
R947 vpwr.n43 vpwr.n40 292.5
R948 vpwr.n45 vpwr.n44 292.5
R949 vpwr.t24 vpwr.t10 287.072
R950 vpwr.t16 vpwr.t8 287.072
R951 vpwr.t12 vpwr.t14 272.274
R952 vpwr.t3 vpwr.t15 254.518
R953 vpwr.t5 vpwr.t18 248.599
R954 vpwr.t15 vpwr.t26 248.599
R955 vpwr.t22 vpwr.t1 244.306
R956 vpwr.n6 vpwr.t31 187.321
R957 vpwr vpwr.t22 186.556
R958 vpwr.n44 vpwr.n43 182.929
R959 vpwr.n7 vpwr.n5 152
R960 vpwr.n42 vpwr.n41 148.689
R961 vpwr.n14 vpwr.t30 126.127
R962 vpwr.n39 vpwr.t27 119.608
R963 vpwr.n58 vpwr.t17 93.81
R964 vpwr.n6 vpwr.n1 73.2067
R965 vpwr.n43 vpwr.t19 68.0124
R966 vpwr.n58 vpwr.t9 63.3219
R967 vpwr.n39 vpwr.t6 63.3219
R968 vpwr.n41 vpwr.t25 61.9158
R969 vpwr.n31 vpwr.t2 41.5552
R970 vpwr.n31 vpwr.t23 41.5552
R971 vpwr.n71 vpwr.n70 34.6358
R972 vpwr.n64 vpwr.n34 34.6358
R973 vpwr.n65 vpwr.n64 34.6358
R974 vpwr.n66 vpwr.n65 34.6358
R975 vpwr.n60 vpwr.n57 34.6358
R976 vpwr.n51 vpwr.n37 34.6358
R977 vpwr.n55 vpwr.n37 34.6358
R978 vpwr.n66 vpwr.n32 32.377
R979 vpwr.n56 vpwr.n55 32.0005
R980 vpwr.n41 vpwr.t11 30.239
R981 vpwr.n50 vpwr.n49 30.1181
R982 vpwr.n44 vpwr.t29 29.316
R983 vpwr.n72 vpwr.n71 22.9652
R984 vpwr.n51 vpwr.n50 20.3299
R985 vpwr.n70 vpwr.n32 18.0711
R986 vpwr vpwr.n4 14.0185
R987 vpwr.n45 vpwr.n42 13.9946
R988 vpwr.n49 vpwr.n40 12.8758
R989 vpwr.n57 vpwr.n56 9.41227
R990 vpwr.n11 vpwr.n10 9.3005
R991 vpwr.n8 vpwr.n2 9.3005
R992 vpwr.n8 vpwr.n7 9.3005
R993 vpwr.n7 vpwr.n6 9.15991
R994 vpwr.n15 vpwr.n14 7.02651
R995 vpwr.n59 vpwr.n34 6.02403
R996 vpwr.n46 vpwr.n45 5.00414
R997 vpwr.n4 vpwr 4.7293
R998 vpwr.n9 vpwr.n0 4.6505
R999 vpwr.n18 vpwr.n17 4.6505
R1000 vpwr.n47 vpwr.n46 4.6505
R1001 vpwr.n49 vpwr.n48 4.6505
R1002 vpwr.n50 vpwr.n38 4.6505
R1003 vpwr.n52 vpwr.n51 4.6505
R1004 vpwr.n53 vpwr.n37 4.6505
R1005 vpwr.n55 vpwr.n54 4.6505
R1006 vpwr.n56 vpwr.n36 4.6505
R1007 vpwr.n57 vpwr.n35 4.6505
R1008 vpwr.n61 vpwr.n60 4.6505
R1009 vpwr.n62 vpwr.n34 4.6505
R1010 vpwr.n64 vpwr.n63 4.6505
R1011 vpwr.n65 vpwr.n33 4.6505
R1012 vpwr.n67 vpwr.n66 4.6505
R1013 vpwr.n68 vpwr.n32 4.6505
R1014 vpwr.n70 vpwr.n69 4.6505
R1015 vpwr.n71 vpwr.n30 4.6505
R1016 vpwr.n4 vpwr 4.53383
R1017 vpwr.n46 vpwr.n40 4.07323
R1018 vpwr.n73 vpwr.n72 3.93272
R1019 vpwr.n60 vpwr.n59 3.76521
R1020 vpwr.n5 vpwr 3.11401
R1021 vpwr.n17 vpwr.n15 3.0725
R1022 vpwr.n27 vpwr.n26 2.91783
R1023 vpwr.n28 vpwr 2.44425
R1024 vpwr.n12 vpwr 2.36657
R1025 vpwr.n5 vpwr.n1 1.55726
R1026 vpwr.n10 vpwr.n9 1.55726
R1027 vpwr.n8 vpwr.n1 1.38428
R1028 vpwr.n9 vpwr.n8 1.38428
R1029 vpwr.n10 vpwr 1.38428
R1030 vpwr.n17 vpwr.n16 1.2805
R1031 vpwr.n77 vpwr.n76 0.711611
R1032 vpwr.n12 vpwr 0.580857
R1033 vpwr.n29 vpwr.n28 0.5255
R1034 vpwr.n75 vpwr 0.223
R1035 vpwr.n3 vpwr 0.196446
R1036 vpwr.n20 vpwr 0.171696
R1037 vpwr.n47 vpwr.n42 0.144332
R1038 vpwr.n73 vpwr.n30 0.138831
R1039 vpwr.n48 vpwr.n47 0.120292
R1040 vpwr.n48 vpwr.n38 0.120292
R1041 vpwr.n52 vpwr.n38 0.120292
R1042 vpwr.n53 vpwr.n52 0.120292
R1043 vpwr.n54 vpwr.n53 0.120292
R1044 vpwr.n54 vpwr.n36 0.120292
R1045 vpwr.n36 vpwr.n35 0.120292
R1046 vpwr.n61 vpwr.n35 0.120292
R1047 vpwr.n62 vpwr.n61 0.120292
R1048 vpwr.n63 vpwr.n62 0.120292
R1049 vpwr.n63 vpwr.n33 0.120292
R1050 vpwr.n67 vpwr.n33 0.120292
R1051 vpwr.n68 vpwr.n67 0.120292
R1052 vpwr.n69 vpwr.n68 0.120292
R1053 vpwr.n69 vpwr.n30 0.120292
R1054 vpwr.n74 vpwr.n73 0.107496
R1055 vpwr.n20 vpwr.n19 0.0901739
R1056 vpwr vpwr.n83 0.0634013
R1057 vpwr.n27 vpwr 0.063
R1058 vpwr.n21 vpwr.n20 0.0500874
R1059 vpwr.n13 vpwr.n12 0.0466957
R1060 vpwr.n24 vpwr.n23 0.0435328
R1061 vpwr.n83 vpwr.n29 0.039096
R1062 vpwr.n18 vpwr.n13 0.0331087
R1063 vpwr.n83 vpwr.n82 0.0287348
R1064 vpwr.n3 vpwr.n2 0.02675
R1065 vpwr vpwr.n11 0.0255
R1066 vpwr.n22 vpwr.n21 0.0213989
R1067 vpwr.n78 vpwr.n75 0.0207266
R1068 vpwr.n26 vpwr.n25 0.018111
R1069 vpwr.n74 vpwr 0.0174271
R1070 vpwr vpwr.n74 0.01675
R1071 vpwr.n19 vpwr.n18 0.014087
R1072 vpwr.n24 vpwr.n22 0.0127951
R1073 vpwr.n11 vpwr.n0 0.01175
R1074 vpwr.n2 vpwr.n0 0.0105
R1075 vpwr.n81 vpwr.n80 0.009875
R1076 vpwr vpwr.n3 0.00725676
R1077 vpwr.n23 vpwr 0.00459836
R1078 vpwr.n79 vpwr.n78 0.00412592
R1079 vpwr.n80 vpwr.n79 0.003625
R1080 vpwr.n82 vpwr.n81 0.00196888
R1081 vpwr.n26 vpwr.n24 0.0016109
R1082 vpwr.n78 vpwr.n77 0.00154933
R1083 vpwr.n28 vpwr.n27 0.000500433
R1084 vtd.n7 vtd.t29 64.6821
R1085 vtd.n8 vtd.t27 64.3461
R1086 vtd.n4 vtd.t24 63.6317
R1087 vtd.n9 vtd.t26 63.6292
R1088 vtd.n8 vtd.t28 63.6292
R1089 vtd.n17 vtd.t8 63.6292
R1090 vtd.n2 vtd.t6 63.6292
R1091 vtd.n18 vtd.t14 63.6292
R1092 vtd.n1 vtd.t10 63.6292
R1093 vtd.n19 vtd.t12 63.6292
R1094 vtd.n0 vtd.t2 63.6292
R1095 vtd.n6 vtd.t4 63.6292
R1096 vtd.n3 vtd.t0 63.6275
R1097 vtd.n13 vtd.t20 18.2948
R1098 vtd.n10 vtd.t17 18.1899
R1099 vtd.n10 vtd.t21 17.4187
R1100 vtd.n13 vtd.t16 17.4177
R1101 vtd.n11 vtd.t18 17.4156
R1102 vtd.n14 vtd.t23 17.4136
R1103 vtd.n12 vtd.t22 17.4125
R1104 vtd.n15 vtd.t19 17.4115
R1105 vtd.n3 vtd.t1 14.3559
R1106 vtd.n17 vtd.t9 14.3555
R1107 vtd.n2 vtd.t15 14.283
R1108 vtd.n2 vtd.t7 14.283
R1109 vtd.n1 vtd.t13 14.283
R1110 vtd.n1 vtd.t11 14.283
R1111 vtd.n0 vtd.t5 14.283
R1112 vtd.n0 vtd.t3 14.283
R1113 vtd.n7 vtd.t25 13.7801
R1114 vtd.n16 vtd.n15 2.14635
R1115 vtd.n3 vtd.n16 1.54335
R1116 vtd vtd.n20 1.22372
R1117 vtd.n16 vtd.n12 1.09526
R1118 vtd.n20 vtd.n3 0.981002
R1119 vtd.n15 vtd.n14 0.8755
R1120 vtd.n14 vtd.n13 0.8755
R1121 vtd.n5 vtd.n7 0.832184
R1122 vtd.n11 vtd.n10 0.769433
R1123 vtd.n12 vtd.n11 0.769356
R1124 vtd.n9 vtd.n8 0.717388
R1125 vtd.n4 vtd.n9 0.708453
R1126 vtd.n20 vtd.n5 0.438348
R1127 vtd.n3 vtd.n6 0.140567
R1128 vtd.n18 vtd.n2 0.140142
R1129 vtd.n19 vtd.n1 0.140142
R1130 vtd.n6 vtd.n0 0.140142
R1131 vtd.n0 vtd.n19 0.134875
R1132 vtd.n1 vtd.n18 0.134875
R1133 vtd.n2 vtd.n17 0.134875
R1134 vtd.n5 vtd.n4 0.114328
R1135 vts.n5 vts.t5 1023.62
R1136 vts.n0 vts.n5 641.967
R1137 vts.t1 vts.t12 333.303
R1138 vts.n0 vts.t1 237.054
R1139 vts.t12 vts.t10 229.925
R1140 vts.t23 vts.t8 229.925
R1141 vts.t21 vts.t19 229.925
R1142 vts.t19 vts.t17 229.925
R1143 vts.t17 vts.t15 229.925
R1144 vts.n5 vts.t23 130.113
R1145 vts.n5 vts.t21 99.8157
R1146 vts.n15 vts.t4 63.6292
R1147 vts.n18 vts.t0 63.6292
R1148 vts.n7 vts.t31 27.6073
R1149 vts.n12 vts.t32 27.1628
R1150 vts.n11 vts.t25 26.7019
R1151 vts.n6 vts.t26 26.4053
R1152 vts.n6 vts.t34 26.2229
R1153 vts.n10 vts.t30 25.2012
R1154 vts.n8 vts.t33 25.2012
R1155 vts.n13 vts.t27 24.699
R1156 vts.n9 vts.t28 24.699
R1157 vts.n14 vts.t29 24.1526
R1158 vts.n0 vts.t14 16.8006
R1159 vts.n16 vts.t6 14.4639
R1160 vts.n17 vts.t3 14.4362
R1161 vts.n19 vts.t2 14.4313
R1162 vts.n15 vts.t7 14.3697
R1163 vts.n1 vts.t13 14.283
R1164 vts.n1 vts.t11 14.283
R1165 vts.n2 vts.t22 14.283
R1166 vts.n2 vts.t20 14.283
R1167 vts.n3 vts.t18 14.283
R1168 vts.n3 vts.t16 14.283
R1169 vts.n4 vts.t9 14.283
R1170 vts.n4 vts.t24 14.283
R1171 vts vts.n14 2.98635
R1172 vts.n11 vts.n10 2.30564
R1173 vts.n7 vts.n6 2.30482
R1174 vts.n9 vts.n8 2.27981
R1175 vts.n13 vts.n12 2.24388
R1176 vts vts.n20 0.8255
R1177 vts.n12 vts.n11 0.680761
R1178 vts.n10 vts.n9 0.680308
R1179 vts.n14 vts.n13 0.680308
R1180 vts.n1 vts.n4 0.65792
R1181 vts.n4 vts.n2 0.65792
R1182 vts.n2 vts.n3 0.6455
R1183 vts.n8 vts.n7 0.604164
R1184 vts.n3 vts.n16 0.462781
R1185 vts.n17 vts.n1 0.452971
R1186 vts.n0 vts.n19 0.0947919
R1187 vts.n16 vts.n15 0.0741592
R1188 vts.n18 vts.n17 0.0682354
R1189 vts.n20 vts.n0 0.0679811
R1190 vts.n19 vts.n18 0.0634447
R1191 buffer_0.b.n0 buffer_0.b.t11 40.2461
R1192 buffer_0.b.n2 buffer_0.b.t10 40.2461
R1193 buffer_0.b buffer_0.b.t9 39.5317
R1194 buffer_0.b.n1 buffer_0.b.t16 39.5292
R1195 buffer_0.b.n1 buffer_0.b.t18 39.5292
R1196 buffer_0.b.n0 buffer_0.b.t13 39.5292
R1197 buffer_0.b.n0 buffer_0.b.t14 39.5292
R1198 buffer_0.b.n3 buffer_0.b.t12 39.5292
R1199 buffer_0.b.n3 buffer_0.b.t19 39.5292
R1200 buffer_0.b.n2 buffer_0.b.t17 39.5292
R1201 buffer_0.b.n2 buffer_0.b.t15 39.5292
R1202 buffer_0.b.n4 buffer_0.b.t1 17.4005
R1203 buffer_0.b.n4 buffer_0.b.t5 17.4005
R1204 buffer_0.b.n6 buffer_0.b.t8 17.4005
R1205 buffer_0.b.n6 buffer_0.b.t4 17.4005
R1206 buffer_0.b.n7 buffer_0.b.t3 17.4005
R1207 buffer_0.b.n7 buffer_0.b.t7 17.4005
R1208 buffer_0.b.n5 buffer_0.b.t6 17.4005
R1209 buffer_0.b.n5 buffer_0.b.t0 17.4005
R1210 buffer_0.b.n4 buffer_0.b.n5 3.1733
R1211 buffer_0.b.n6 buffer_0.b.n7 2.69321
R1212 buffer_0.b.n5 buffer_0.b.n6 2.68836
R1213 buffer_0.b.t2 buffer_0.b.n4 2.65092
R1214 buffer_0.b.n3 buffer_0.b.n2 2.15117
R1215 buffer_0.b.n1 buffer_0.b.n0 2.15117
R1216 buffer_0.b buffer_0.b.n1 1.49152
R1217 buffer_0.b buffer_0.b.t2 0.968485
R1218 buffer_0.b buffer_0.b.n3 0.961845
R1219 buffer_0.c buffer_0.c.t20 18.4486
R1220 buffer_0.c.n17 buffer_0.c.t5 17.4005
R1221 buffer_0.c.n17 buffer_0.c.t16 17.4005
R1222 buffer_0.c.n15 buffer_0.c.t17 17.4005
R1223 buffer_0.c.n15 buffer_0.c.t7 17.4005
R1224 buffer_0.c.n13 buffer_0.c.t2 17.4005
R1225 buffer_0.c.n13 buffer_0.c.t11 17.4005
R1226 buffer_0.c.n9 buffer_0.c.t4 17.4005
R1227 buffer_0.c.n9 buffer_0.c.t19 17.4005
R1228 buffer_0.c.n7 buffer_0.c.t14 17.4005
R1229 buffer_0.c.n7 buffer_0.c.t6 17.4005
R1230 buffer_0.c.n5 buffer_0.c.t1 17.4005
R1231 buffer_0.c.n5 buffer_0.c.t13 17.4005
R1232 buffer_0.c.n3 buffer_0.c.t10 17.4005
R1233 buffer_0.c.n3 buffer_0.c.t3 17.4005
R1234 buffer_0.c.n1 buffer_0.c.t0 17.4005
R1235 buffer_0.c.n1 buffer_0.c.t18 17.4005
R1236 buffer_0.c.n0 buffer_0.c.t15 17.4005
R1237 buffer_0.c.n0 buffer_0.c.t8 17.4005
R1238 buffer_0.c.n11 buffer_0.c.t12 17.4005
R1239 buffer_0.c.n11 buffer_0.c.t9 17.4005
R1240 buffer_0.c.n2 buffer_0.c.n0 1.87829
R1241 buffer_0.c buffer_0.c.n18 1.52139
R1242 buffer_0.c.n18 buffer_0.c.n17 1.51465
R1243 buffer_0.c.n4 buffer_0.c.n2 1.08383
R1244 buffer_0.c.n6 buffer_0.c.n4 1.08383
R1245 buffer_0.c.n10 buffer_0.c.n8 1.08383
R1246 buffer_0.c.n12 buffer_0.c.n10 1.08383
R1247 buffer_0.c.n14 buffer_0.c.n12 1.08383
R1248 buffer_0.c.n8 buffer_0.c.n6 1.04217
R1249 buffer_0.c.n16 buffer_0.c.n14 1.04217
R1250 buffer_0.c.n6 buffer_0.c.n5 0.776026
R1251 buffer_0.c.n14 buffer_0.c.n13 0.766495
R1252 buffer_0.c.n4 buffer_0.c.n3 0.766495
R1253 buffer_0.c.n16 buffer_0.c.n15 0.766495
R1254 buffer_0.c.n10 buffer_0.c.n9 0.766495
R1255 buffer_0.c.n8 buffer_0.c.n7 0.766495
R1256 buffer_0.c.n2 buffer_0.c.n1 0.766495
R1257 buffer_0.c.n12 buffer_0.c.n11 0.766495
R1258 buffer_0.c.n18 buffer_0.c.n16 0.333833
R1259 ib.n1 ib.t5 38.0465
R1260 ib.n1 ib.t3 37.3602
R1261 ib.n3 ib.t0 18.7313
R1262 ib.n3 ib.t2 17.409
R1263 ib.n0 ib.t4 17.4005
R1264 ib.n0 ib.t1 17.4005
R1265 ib ib.n4 1.76488
R1266 ib.n2 ib.n1 0.239515
R1267 ib.n4 ib.n3 0.0163842
R1268 ib.n2 ib.n0 0.00444823
R1269 ib.n4 ib.n2 0.00358796
R1270 out_sigma.n0 out_sigma.t2 394.808
R1271 out_sigma.n1 out_sigma.t0 250.94
R1272 out_sigma out_sigma.t1 144.601
R1273 out_sigma out_sigma.n0 9.0826
R1274 out_sigma.n1 out_sigma 4.7225
R1275 out_sigma out_sigma.n1 3.35288
R1276 out_sigma.n0 out_sigma 0.727062
R1277 clk.n0 clk.t0 294.557
R1278 clk.n0 clk.t1 211.01
R1279 clk.n2 clk.n0 8.28655
R1280 clk.n3 clk 7.73487
R1281 clk.n3 clk.n2 1.82961
R1282 clk.n1 clk 0.981259
R1283 clk.n2 clk.n1 0.848973
R1284 clk clk.n5 0.385917
R1285 clk.n5 clk.n4 0.03175
R1286 clk.n4 clk.n3 0.00111796
R1287 out.n2 out.t0 8.97158
R1288 out.n2 out.n1 2.56714
R1289 out.n0 out.t2 0.506271
R1290 out.n1 out.n0 0.504061
R1291 out out.n2 0.240344
R1292 out.n0 out.t1 0.0277714
R1293 out.n1 out.t3 0.00303875
C0 sigma-delta_0.x1.D vpwr 0.483f
C1 a_14625_2515# clk 0.274f
C2 sigma-delta_0.x1.D sigma-delta_0.x1.Q 0.0675f
C3 vpwr a_15048_3988# 0.00379f
C4 sensor_0.b ib 2.02e-19
C5 buffer_0.d ib 0.194f
C6 a_16024_5320# a_15546_5320# 0.144f
C7 sigma-delta_0.x1.D a_15359_2757# 6.24e-19
C8 a_14550_5320# out 0.00197f
C9 a_15046_2515# a_14791_2515# 0.0642f
C10 a_6126_29386# out 0.0171f
C11 a_15881_2489# a_16522_3988# 1.28e-20
C12 a_15706_2515# a_15868_2881# 0.00645f
C13 vd a_16854_3988# 0.0174f
C14 out_sigma clk 0.11f
C15 out a_16024_5320# 0.00189f
C16 a_14625_2515# a_14716_3988# 1.47e-19
C17 vpwr a_16060_2515# 0.00312f
C18 sigma-delta_0.x1.Q a_16060_2515# 6.05e-19
C19 a_15237_2515# a_14791_2515# 2.28e-19
C20 vd vpwr 0.00726f
C21 a_14550_5320# vd 0.067f
C22 sigma-delta_0.x1.Q vd 0.0969f
C23 a_6126_29386# vd 0.0189f
C24 buffer_0.a buffer_0.c 3.88f
C25 out_buff a_15214_5320# 5.44e-19
C26 vd a_16024_5320# 0.0626f
C27 a_15712_3988# a_14716_3988# 2.04e-19
C28 vd sensor_0.c 0.804f
C29 buffer_0.d out 0.00472f
C30 out_sigma a_14716_3988# 0.0146f
C31 a_16445_2515# a_15706_2515# 7.05e-19
C32 a_15046_2515# clk 3.09e-19
C33 a_15712_3988# a_17020_5320# 0.00974f
C34 sigma-delta_0.x1.D a_15868_2881# 2.11e-20
C35 a_14625_2515# a_15712_3988# 1.78e-19
C36 buffer_0.c ib 0.0951f
C37 a_14625_2515# out_sigma 0.00153f
C38 vpwr a_14791_2515# 0.607f
C39 sigma-delta_0.x1.Q a_14791_2515# 0.00137f
C40 vd sensor_0.b 0.0693f
C41 vd buffer_0.d 2.79f
C42 a_15237_2515# clk 5.33e-20
C43 a_15706_2515# a_15141_2515# 7.99e-20
C44 a_15048_3988# a_14882_5320# 0.00482f
C45 vpwr a_15881_2489# 0.688f
C46 sensor_0.c sensor_0.a 0.997f
C47 sigma-delta_0.x1.Q a_15881_2489# 0.142f
C48 a_15141_2515# a_15380_3988# 1.22e-19
C49 a_15359_2757# a_14791_2515# 0.186f
C50 vd a_16190_3988# 0.00388f
C51 buffer_0.b buffer_0.d 1.04f
C52 buffer_0.a out_buff 3.96f
C53 a_15712_3988# out_sigma 0.16f
C54 out a_14882_5320# 0.0019f
C55 sigma-delta_0.x1.D a_15249_2881# 5.56e-20
C56 vts sensor_0.c 0.192f
C57 out a_16356_5320# 0.00195f
C58 sensor_0.b sensor_0.a 0.821f
C59 a_16445_2515# sigma-delta_0.x1.D 0.00209f
C60 a_14625_2515# a_15046_2515# 0.0931f
C61 out_buff a_15380_3988# 4.51e-19
C62 vpwr clk 0.729f
C63 out_buff ib 0.0112f
C64 vd a_14882_5320# 0.061f
C65 out buffer_0.c 8.56e-19
C66 a_15712_3988# a_16522_3988# 0.0502f
C67 vd a_16356_5320# 0.0637f
C68 vts sensor_0.b 0.974f
C69 buffer_0.d vts 0.213f
C70 sigma-delta_0.x1.D a_15141_2515# 0.00353f
C71 a_14625_2515# a_15237_2515# 0.00134f
C72 a_15214_5320# a_15380_3988# 0.00473f
C73 a_15359_2757# clk 1.78e-19
C74 a_15881_2489# a_16190_3988# 4.27e-19
C75 a_15403_2515# sigma-delta_0.x1.D 5.41e-20
C76 vd buffer_0.c 0.399f
C77 a_14791_2515# a_15868_2881# 1.46e-19
C78 a_16854_3988# a_17020_5320# 0.00434f
C79 a_16445_2515# vd 0.00317f
C80 out_buff a_15546_5320# 2.84e-19
C81 vpwr a_14716_3988# 0.0038f
C82 a_14550_5320# a_14716_3988# 0.00458f
C83 out_buff a_15048_3988# 0.00101f
C84 buffer_0.b buffer_0.c 1.34f
C85 buffer_0.d clk 0.205f
C86 sigma-delta_0.x1.Q a_17020_5320# 0.00839f
C87 a_15706_2515# a_15815_2515# 0.00742f
C88 a_14625_2515# vpwr 0.772f
C89 a_15214_5320# a_15546_5320# 0.296f
C90 a_14625_2515# sigma-delta_0.x1.Q 9.54e-19
C91 a_15048_3988# a_15214_5320# 0.00473f
C92 a_15712_3988# a_16854_3988# 0.00957f
C93 out_buff out 0.0109f
C94 a_14791_2515# a_15249_2881# 0.0346f
C95 out_sigma a_16854_3988# 7.61e-19
C96 a_14625_2515# a_15359_2757# 0.0701f
C97 buffer_0.a ib 0.0615f
C98 a_16445_2515# a_14791_2515# 2.01e-19
C99 a_15712_3988# vpwr 0.0132f
C100 a_15712_3988# sigma-delta_0.x1.Q 0.414f
C101 out a_15214_5320# 0.00184f
C102 vts buffer_0.c 1.08f
C103 out_sigma a_14550_5320# 6.23e-19
C104 out_sigma vpwr 0.597f
C105 sigma-delta_0.x1.Q out_sigma 0.668f
C106 a_15237_2515# a_15046_2515# 4.61e-19
C107 vd out_buff 3.21f
C108 a_16445_2515# a_15881_2489# 0.107f
C109 a_16688_5320# out 0.00185f
C110 a_15712_3988# a_16024_5320# 0.00827f
C111 a_15141_2515# a_14791_2515# 0.23f
C112 a_15712_3988# a_15359_2757# 7.49e-21
C113 a_16854_3988# a_16522_3988# 0.303f
C114 vd sensor_0.d 0.282f
C115 out_sigma a_15359_2757# 3.73e-19
C116 buffer_0.b out_buff 2.8f
C117 sigma-delta_0.x1.D a_15815_2515# 2.42e-20
C118 vd a_15214_5320# 0.0598f
C119 vpwr a_16522_3988# 0.00266f
C120 a_16688_5320# vd 0.0633f
C121 sigma-delta_0.x1.Q a_16522_3988# 5e-20
C122 sigma-delta_0.x1.D a_15706_2515# 9.45e-19
C123 vpwr a_15046_2515# 0.0861f
C124 a_15380_3988# a_15546_5320# 0.00434f
C125 sigma-delta_0.x1.Q a_15046_2515# 7.58e-20
C126 buffer_0.a out 0.0533f
C127 out_sigma buffer_0.d 0.0399f
C128 a_14716_3988# a_14882_5320# 0.00434f
C129 sensor_0.d sensor_0.a 0.588f
C130 a_15048_3988# a_15380_3988# 0.302f
C131 a_15712_3988# a_16190_3988# 0.357f
C132 out_buff vts 2.36f
C133 a_15141_2515# clk 3.26e-19
C134 a_15237_2515# vpwr 0.00292f
C135 sigma-delta_0.x1.Q a_15237_2515# 1.45e-19
C136 buffer_0.a vd 6.66f
C137 vts sensor_0.d 0.248f
C138 a_15403_2515# clk 1.82e-20
C139 a_15712_3988# a_15868_2881# 5.54e-20
C140 a_15237_2515# a_15359_2757# 3.16e-19
C141 buffer_0.a buffer_0.b 0.126f
C142 a_14625_2515# a_15249_2881# 9.73e-19
C143 a_15706_2515# vd 3.52e-19
C144 sigma-delta_0.x1.Q a_16854_3988# 0.414f
C145 a_16190_3988# a_16522_3988# 0.312f
C146 out_buff clk 0.0713f
C147 a_15712_3988# a_16356_5320# 0.00631f
C148 vd a_15380_3988# 0.00209f
C149 a_16445_2515# a_14625_2515# 4.71e-20
C150 sigma-delta_0.x1.D a_15048_3988# 2.56e-20
C151 vd ib 0.0605f
C152 a_15815_2515# a_14791_2515# 2.36e-20
C153 sigma-delta_0.x1.Q vpwr 0.186f
C154 out a_15546_5320# 0.00187f
C155 a_14625_2515# a_15141_2515# 0.115f
C156 buffer_0.b ib 0.0167f
C157 out_sigma buffer_0.c 0.00107f
C158 vpwr a_15359_2757# 0.378f
C159 a_16445_2515# a_15712_3988# 0.00366f
C160 sigma-delta_0.x1.Q a_15359_2757# 0.00111f
C161 buffer_0.a vts 0.658f
C162 a_16445_2515# out_sigma 0.0691f
C163 a_15706_2515# a_14791_2515# 0.125f
C164 a_16522_3988# a_16356_5320# 0.00509f
C165 out_buff a_14716_3988# 0.306f
C166 vd a_15546_5320# 0.0619f
C167 sigma-delta_0.x1.D a_16060_2515# 4.54e-20
C168 sigma-delta_0.x1.D vd 0.908f
C169 a_15712_3988# a_15141_2515# 2.02e-20
C170 a_15706_2515# a_15881_2489# 0.251f
C171 vd a_15048_3988# 0.00206f
C172 a_15141_2515# out_sigma 7.05e-19
C173 a_15815_2515# clk 1.1e-20
C174 vts ib 0.723f
C175 a_16445_2515# a_16522_3988# 1.4e-19
C176 vd out 0.145p
C177 vpwr a_16190_3988# 0.00384f
C178 sigma-delta_0.x1.Q a_16190_3988# 1.87e-20
C179 sensor_0.b sensor_0.c 0.55f
C180 a_15712_3988# out_buff 0.00915f
C181 a_16688_5320# a_17020_5320# 0.299f
C182 buffer_0.b out 0.0634f
C183 out_sigma out_buff 0.552f
C184 a_15706_2515# clk 6.46e-20
C185 a_16024_5320# a_16190_3988# 0.00473f
C186 sigma-delta_0.x1.D a_14791_2515# 0.229f
C187 vpwr a_15868_2881# 9.63e-19
C188 a_14791_2515# a_15048_3988# 1.82e-19
C189 sigma-delta_0.x1.Q a_15868_2881# 4.53e-20
C190 a_15141_2515# a_15046_2515# 0.0498f
C191 sigma-delta_0.x1.D a_15881_2489# 0.004f
C192 a_14550_5320# a_14882_5320# 0.296f
C193 a_15359_2757# a_15868_2881# 2.6e-19
C194 buffer_0.b vd 6.37f
C195 a_16688_5320# a_15712_3988# 0.00557f
C196 a_14625_2515# a_15815_2515# 2.56e-19
C197 a_15141_2515# a_15237_2515# 0.0138f
C198 vts out 0.00336f
C199 a_16024_5320# a_16356_5320# 0.3f
C200 vd sensor_0.a 2.92f
C201 vpwr a_15249_2881# 0.156f
C202 sigma-delta_0.x1.Q a_15249_2881# 3.66e-19
C203 vd a_14791_2515# 1.08e-19
C204 a_16445_2515# vpwr 0.2f
C205 sigma-delta_0.x1.D clk 0.00993f
C206 a_14625_2515# a_15706_2515# 0.102f
C207 a_16445_2515# sigma-delta_0.x1.Q 0.226f
C208 a_15712_3988# a_15815_2515# 1.36e-20
C209 a_15881_2489# a_16060_2515# 0.0074f
C210 a_16688_5320# a_16522_3988# 0.00482f
C211 vd a_15881_2489# 0.00172f
C212 vd vts 1.62f
C213 a_15359_2757# a_15249_2881# 0.0977f
C214 buffer_0.a out_sigma 0.0172f
C215 a_15141_2515# vpwr 0.363f
C216 sigma-delta_0.x1.Q a_15141_2515# 8.11e-19
C217 buffer_0.b vts 2.94f
C218 a_15712_3988# a_15706_2515# 0.0011f
C219 a_16190_3988# a_16356_5320# 0.00536f
C220 a_15403_2515# vpwr 0.00407f
C221 a_15706_2515# out_sigma 6.85e-19
C222 a_15403_2515# sigma-delta_0.x1.Q 9.75e-20
C223 a_15712_3988# a_15380_3988# 0.298f
C224 a_15141_2515# a_15359_2757# 0.21f
C225 sigma-delta_0.x1.D a_14716_3988# 2.07e-19
C226 out_sigma a_15380_3988# 0.0148f
C227 buffer_0.d buffer_0.c 1.32f
C228 a_15048_3988# a_14716_3988# 0.296f
C229 a_16060_2515# clk 6.32e-21
C230 vts sensor_0.a 0.543f
C231 a_15881_2489# a_14791_2515# 0.0426f
C232 a_15403_2515# a_15359_2757# 3.69e-19
C233 out_buff vpwr 0.0083f
C234 a_14550_5320# out_buff 0.0535f
C235 a_14625_2515# sigma-delta_0.x1.D 0.195f
C236 a_14625_2515# a_15048_3988# 1.92e-19
C237 a_16688_5320# a_16854_3988# 0.00473f
C238 out_buff a_16024_5320# 3.49e-20
C239 out a_17020_5320# 0.00192f
C240 a_15712_3988# a_15546_5320# 0.00466f
C241 sigma-delta_0.x1.D a_15712_3988# 0.339f
C242 a_16688_5320# sigma-delta_0.x1.Q 0.0032f
C243 a_15712_3988# a_15048_3988# 4.38e-19
C244 vd a_14716_3988# 0.0021f
C245 sigma-delta_0.x1.D out_sigma 0.294f
C246 a_14791_2515# clk 0.00241f
C247 sensor_0.c sensor_0.d 0.492f
C248 out_sigma a_15048_3988# 0.0146f
C249 vd a_17020_5320# 0.201f
C250 buffer_0.d out_buff 40f
C251 a_14625_2515# vd 1.72e-20
C252 a_15881_2489# clk 2.68e-20
C253 a_15712_3988# out 0.18f
C254 out_sigma out 5.44f
C255 sensor_0.b sensor_0.d 0.0152f
C256 out_buff a_16190_3988# 9.87e-22
C257 a_15815_2515# vpwr 7.93e-19
C258 sigma-delta_0.x1.Q a_15815_2515# 1.47e-19
C259 a_15712_3988# vd 0.75f
C260 sigma-delta_0.x1.D a_15046_2515# 0.164f
C261 a_15815_2515# a_15359_2757# 4.2e-19
C262 out_sigma vd 1.88f
C263 a_15706_2515# vpwr 0.524f
C264 a_15706_2515# sigma-delta_0.x1.Q 0.00593f
C265 a_15141_2515# a_15249_2881# 0.0572f
C266 a_14625_2515# a_14791_2515# 0.906f
C267 vpwr a_15380_3988# 0.00397f
C268 sigma-delta_0.x1.Q a_15380_3988# 1.43e-21
C269 buffer_0.b out_sigma 0.017f
C270 out_buff a_14882_5320# 0.0014f
C271 sigma-delta_0.x1.D a_15237_2515# 8.22e-19
C272 a_14625_2515# a_15881_2489# 0.0436f
C273 a_15706_2515# a_15359_2757# 0.0512f
C274 vd a_16522_3988# 0.00558f
C275 a_15359_2757# a_15380_3988# 7.2e-20
C276 a_15214_5320# a_14882_5320# 0.303f
C277 a_15712_3988# a_14791_2515# 4.13e-19
C278 buffer_0.a buffer_0.d 2.4f
C279 sensor_0.c ib 0.00238f
C280 out_sigma a_14791_2515# 0.0011f
C281 out_buff buffer_0.c 2.02f
C282 sigma-delta_0.x1.D a_16854_3988# 2.69e-19
C283 a_16688_5320# a_16356_5320# 0.307f
C284 a_15403_2515# a_15141_2515# 0.00171f
C285 a_15712_3988# a_15881_2489# 0.00381f
C286 out_sigma a_15881_2489# 0.00735f
C287 out_sigma vts 0.0608f
C288 clk gnd 3.43f
C289 ib gnd 6.69f
C290 out gnd 59.7f
C291 vpwr gnd 7.16f
C292 vd gnd 77.8f
C293 a_16060_2515# gnd 0.00223f
C294 a_15815_2515# gnd 9.68e-19
C295 a_15403_2515# gnd 0.00579f
C296 a_15237_2515# gnd 0.00863f
C297 a_15249_2881# gnd 0.00469f
C298 a_15046_2515# gnd 0.08f
C299 a_16445_2515# gnd 0.213f
C300 a_15706_2515# gnd 0.275f
C301 a_15881_2489# gnd 0.74f
C302 a_15141_2515# gnd 0.281f
C303 a_15359_2757# gnd 0.194f
C304 a_14791_2515# gnd 0.332f
C305 sigma-delta_0.x1.D gnd 2.56f
C306 a_14625_2515# gnd 0.7f
C307 sigma-delta_0.x1.Q gnd 1.09f
C308 a_17020_5320# gnd 0.557f
C309 a_16854_3988# gnd 0.348f
C310 a_16688_5320# gnd 0.388f
C311 a_16522_3988# gnd 0.356f
C312 a_16356_5320# gnd 0.392f
C313 a_16190_3988# gnd 0.357f
C314 a_16024_5320# gnd 0.447f
C315 a_15712_3988# gnd 69.7f
C316 a_15546_5320# gnd 0.449f
C317 a_15380_3988# gnd 0.365f
C318 a_15214_5320# gnd 0.387f
C319 a_15048_3988# gnd 0.364f
C320 a_14882_5320# gnd 0.39f
C321 a_14716_3988# gnd 0.366f
C322 buffer_0.c gnd 2.18f
C323 sensor_0.b gnd 16.7f
C324 sensor_0.c gnd 0.658f
C325 sensor_0.a gnd 5.59f
C326 sensor_0.d gnd 0.293f
C327 a_14550_5320# gnd 0.587f
C328 out_buff gnd 15.1f
C329 buffer_0.d gnd 27.7f
C330 buffer_0.b gnd 4.08f
C331 buffer_0.a gnd 5.13f
C332 out_sigma gnd 15.5f
C333 a_6126_29386# gnd 0.593f
C334 vts gnd 22.4f
C335 out.t0 gnd 0.00791f
C336 out.t3 gnd 13.1f
C337 out.t2 gnd 29f
C338 out.t1 gnd 19.9f
C339 out.n0 gnd 10.6f
C340 out.n1 gnd 16.3f
C341 out.n2 gnd 61.5f
C342 out_sigma.t0 gnd 0.00942f
C343 out_sigma.t2 gnd 0.0205f
C344 out_sigma.n0 gnd 1.8f
C345 out_sigma.n1 gnd 0.155f
C346 out_sigma.t1 gnd 0.00695f
C347 buffer_0.c.t15 gnd 0.0162f
C348 buffer_0.c.t8 gnd 0.0162f
C349 buffer_0.c.n0 gnd 0.356f
C350 buffer_0.c.t0 gnd 0.0162f
C351 buffer_0.c.t18 gnd 0.0162f
C352 buffer_0.c.n1 gnd 0.258f
C353 buffer_0.c.n2 gnd 0.326f
C354 buffer_0.c.t10 gnd 0.0162f
C355 buffer_0.c.t3 gnd 0.0162f
C356 buffer_0.c.n3 gnd 0.258f
C357 buffer_0.c.n4 gnd 0.25f
C358 buffer_0.c.t1 gnd 0.0162f
C359 buffer_0.c.t13 gnd 0.0162f
C360 buffer_0.c.n5 gnd 0.257f
C361 buffer_0.c.n6 gnd 0.249f
C362 buffer_0.c.t14 gnd 0.0162f
C363 buffer_0.c.t6 gnd 0.0162f
C364 buffer_0.c.n7 gnd 0.258f
C365 buffer_0.c.n8 gnd 0.247f
C366 buffer_0.c.t4 gnd 0.0162f
C367 buffer_0.c.t19 gnd 0.0162f
C368 buffer_0.c.n9 gnd 0.258f
C369 buffer_0.c.n10 gnd 0.25f
C370 buffer_0.c.t12 gnd 0.0162f
C371 buffer_0.c.t9 gnd 0.0162f
C372 buffer_0.c.n11 gnd 0.259f
C373 buffer_0.c.n12 gnd 0.25f
C374 buffer_0.c.t2 gnd 0.0162f
C375 buffer_0.c.t11 gnd 0.0162f
C376 buffer_0.c.n13 gnd 0.258f
C377 buffer_0.c.n14 gnd 0.247f
C378 buffer_0.c.t17 gnd 0.0162f
C379 buffer_0.c.t7 gnd 0.0162f
C380 buffer_0.c.n15 gnd 0.258f
C381 buffer_0.c.n16 gnd 0.187f
C382 buffer_0.c.t5 gnd 0.0162f
C383 buffer_0.c.t16 gnd 0.0162f
C384 buffer_0.c.n17 gnd 0.333f
C385 buffer_0.c.n18 gnd 0.298f
C386 buffer_0.c.t20 gnd 0.0328f
C387 buffer_0.b.n0 gnd 0.787f
C388 buffer_0.b.n1 gnd 0.539f
C389 buffer_0.b.n2 gnd 0.787f
C390 buffer_0.b.n3 gnd 0.619f
C391 buffer_0.b.n4 gnd 0.789f
C392 buffer_0.b.n5 gnd 0.719f
C393 buffer_0.b.n6 gnd 0.798f
C394 buffer_0.b.t10 gnd 0.465f
C395 buffer_0.b.t15 gnd 0.46f
C396 buffer_0.b.t17 gnd 0.46f
C397 buffer_0.b.t19 gnd 0.46f
C398 buffer_0.b.t12 gnd 0.46f
C399 buffer_0.b.t9 gnd 0.46f
C400 buffer_0.b.t16 gnd 0.46f
C401 buffer_0.b.t18 gnd 0.46f
C402 buffer_0.b.t13 gnd 0.46f
C403 buffer_0.b.t14 gnd 0.46f
C404 buffer_0.b.t11 gnd 0.465f
C405 buffer_0.b.t1 gnd 0.0187f
C406 buffer_0.b.t5 gnd 0.0187f
C407 buffer_0.b.t8 gnd 0.0187f
C408 buffer_0.b.t4 gnd 0.0187f
C409 buffer_0.b.t3 gnd 0.0187f
C410 buffer_0.b.t7 gnd 0.0187f
C411 buffer_0.b.n7 gnd 0.505f
C412 buffer_0.b.t6 gnd 0.0187f
C413 buffer_0.b.t0 gnd 0.0187f
C414 buffer_0.b.t2 gnd 0.607f
C415 vts.n0 gnd 1.22f
C416 vts.n1 gnd 0.126f
C417 vts.n2 gnd 0.14f
C418 vts.n3 gnd 0.127f
C419 vts.n4 gnd 0.14f
C420 vts.n5 gnd 0.835f
C421 vts.t26 gnd 0.098f
C422 vts.t34 gnd 0.0974f
C423 vts.n6 gnd 0.153f
C424 vts.t31 gnd 0.0998f
C425 vts.n7 gnd 0.0925f
C426 vts.t33 gnd 0.0955f
C427 vts.n8 gnd 0.0994f
C428 vts.t28 gnd 0.0945f
C429 vts.n9 gnd 0.0996f
C430 vts.t30 gnd 0.0955f
C431 vts.n10 gnd 0.097f
C432 vts.t25 gnd 0.0983f
C433 vts.n11 gnd 0.0944f
C434 vts.t32 gnd 0.0991f
C435 vts.n12 gnd 0.094f
C436 vts.t27 gnd 0.0945f
C437 vts.n13 gnd 0.0994f
C438 vts.t29 gnd 0.0933f
C439 vts.n14 gnd 0.141f
C440 vts.t0 gnd 0.174f
C441 vts.t13 gnd 0.00994f
C442 vts.t11 gnd 0.00994f
C443 vts.t22 gnd 0.00994f
C444 vts.t20 gnd 0.00994f
C445 vts.t18 gnd 0.00994f
C446 vts.t16 gnd 0.00994f
C447 vts.t6 gnd 0.0107f
C448 vts.t4 gnd 0.174f
C449 vts.t7 gnd 0.0105f
C450 vts.n15 gnd 0.208f
C451 vts.n16 gnd 0.119f
C452 vts.t9 gnd 0.00994f
C453 vts.t24 gnd 0.00994f
C454 vts.t3 gnd 0.0106f
C455 vts.n17 gnd 0.119f
C456 vts.n18 gnd 0.112f
C457 vts.t2 gnd 0.0106f
C458 vts.n19 gnd 0.0951f
C459 vts.t10 gnd 0.471f
C460 vts.t12 gnd 0.577f
C461 vts.t1 gnd 0.585f
C462 vts.t5 gnd 1.07f
C463 vts.t8 gnd 0.471f
C464 vts.t23 gnd 0.369f
C465 vts.t15 gnd 0.583f
C466 vts.t17 gnd 0.471f
C467 vts.t19 gnd 0.471f
C468 vts.t21 gnd 0.338f
C469 vts.t14 gnd 0.0656f
C470 vts.n20 gnd 0.06f
C471 vtd.n0 gnd 0.548f
C472 vtd.n1 gnd 0.548f
C473 vtd.n2 gnd 0.548f
C474 vtd.n3 gnd 0.963f
C475 vtd.n4 gnd 0.175f
C476 vtd.n5 gnd 0.236f
C477 vtd.n6 gnd 0.323f
C478 vtd.t25 gnd 2.08f
C479 vtd.t29 gnd 0.404f
C480 vtd.n7 gnd 1.27f
C481 vtd.t27 gnd 0.403f
C482 vtd.t28 gnd 0.401f
C483 vtd.n8 gnd 0.398f
C484 vtd.t26 gnd 0.401f
C485 vtd.n9 gnd 0.205f
C486 vtd.t24 gnd 0.401f
C487 vtd.t17 gnd 0.0205f
C488 vtd.t21 gnd 0.0115f
C489 vtd.n10 gnd 0.439f
C490 vtd.t18 gnd 0.0115f
C491 vtd.n11 gnd 0.236f
C492 vtd.t22 gnd 0.0115f
C493 vtd.n12 gnd 0.248f
C494 vtd.t19 gnd 0.0115f
C495 vtd.t16 gnd 0.0115f
C496 vtd.t20 gnd 0.0206f
C497 vtd.n13 gnd 0.4f
C498 vtd.t23 gnd 0.0115f
C499 vtd.n14 gnd 0.22f
C500 vtd.n15 gnd 0.324f
C501 vtd.n16 gnd 0.453f
C502 vtd.t1 gnd 0.024f
C503 vtd.t0 gnd 0.401f
C504 vtd.t4 gnd 0.401f
C505 vtd.t5 gnd 0.0229f
C506 vtd.t3 gnd 0.0229f
C507 vtd.t2 gnd 0.401f
C508 vtd.t12 gnd 0.401f
C509 vtd.t13 gnd 0.0229f
C510 vtd.t11 gnd 0.0229f
C511 vtd.t10 gnd 0.401f
C512 vtd.t14 gnd 0.401f
C513 vtd.t15 gnd 0.0229f
C514 vtd.t7 gnd 0.0229f
C515 vtd.t6 gnd 0.401f
C516 vtd.t8 gnd 0.401f
C517 vtd.t9 gnd 0.0239f
C518 vtd.n17 gnd 0.532f
C519 vtd.n18 gnd 0.341f
C520 vtd.n19 gnd 0.341f
C521 vtd.n20 gnd 0.626f
C522 sensor_0.a.n0 gnd 0.396f
C523 sensor_0.a.n1 gnd 0.413f
C524 sensor_0.a.t15 gnd 0.277f
C525 sensor_0.a.t14 gnd 0.276f
C526 sensor_0.a.n2 gnd 0.293f
C527 sensor_0.a.t12 gnd 0.276f
C528 sensor_0.a.n3 gnd 0.15f
C529 sensor_0.a.t13 gnd 0.276f
C530 sensor_0.a.n4 gnd 0.148f
C531 sensor_0.a.t1 gnd 0.0159f
C532 sensor_0.a.t0 gnd 0.276f
C533 sensor_0.a.t2 gnd 0.276f
C534 sensor_0.a.t3 gnd 0.0177f
C535 sensor_0.a.t11 gnd 0.0141f
C536 sensor_0.a.t8 gnd 0.00791f
C537 sensor_0.a.n5 gnd 0.277f
C538 sensor_0.a.t7 gnd 0.00792f
C539 sensor_0.a.n6 gnd 0.152f
C540 sensor_0.a.t4 gnd 0.00792f
C541 sensor_0.a.n7 gnd 0.19f
C542 sensor_0.a.t6 gnd 0.0141f
C543 sensor_0.a.t10 gnd 0.00791f
C544 sensor_0.a.n8 gnd 0.276f
C545 sensor_0.a.t5 gnd 0.0079f
C546 sensor_0.a.n9 gnd 0.154f
C547 sensor_0.a.t9 gnd 0.00792f
C548 sensor_0.a.n10 gnd 0.19f
C549 sensor_0.a.n11 gnd 0.384f
C550 sensor_0.b.t19 gnd 0.0077f
C551 sensor_0.b.t1 gnd 0.0077f
C552 sensor_0.b.n0 gnd 0.0683f
C553 sensor_0.b.t0 gnd 0.0077f
C554 sensor_0.b.t18 gnd 0.0077f
C555 sensor_0.b.n1 gnd 0.0506f
C556 sensor_0.b.n2 gnd 0.162f
C557 sensor_0.b.t5 gnd 0.00651f
C558 sensor_0.b.t13 gnd 0.00386f
C559 sensor_0.b.n3 gnd 0.139f
C560 sensor_0.b.t7 gnd 0.00385f
C561 sensor_0.b.n4 gnd 0.0928f
C562 sensor_0.b.t15 gnd 0.00385f
C563 sensor_0.b.n5 gnd 0.137f
C564 sensor_0.b.n6 gnd 0.202f
C565 sensor_0.b.t4 gnd 0.134f
C566 sensor_0.b.t12 gnd 0.127f
C567 sensor_0.b.t6 gnd 0.127f
C568 sensor_0.b.t14 gnd 0.0845f
C569 sensor_0.b.t32 gnd 0.134f
C570 sensor_0.b.t24 gnd 0.127f
C571 sensor_0.b.t31 gnd 0.127f
C572 sensor_0.b.t23 gnd 0.0845f
C573 sensor_0.b.t26 gnd 0.134f
C574 sensor_0.b.t34 gnd 0.127f
C575 sensor_0.b.t21 gnd 0.127f
C576 sensor_0.b.t29 gnd 0.0845f
C577 sensor_0.b.t20 gnd 0.134f
C578 sensor_0.b.t27 gnd 0.127f
C579 sensor_0.b.t28 gnd 0.127f
C580 sensor_0.b.t35 gnd 0.0845f
C581 sensor_0.b.t30 gnd 0.134f
C582 sensor_0.b.t22 gnd 0.127f
C583 sensor_0.b.t33 gnd 0.127f
C584 sensor_0.b.t25 gnd 0.0856f
C585 sensor_0.b.n7 gnd 0.119f
C586 sensor_0.b.n8 gnd 0.0626f
C587 sensor_0.b.n9 gnd 0.0626f
C588 sensor_0.b.n10 gnd 0.0626f
C589 sensor_0.b.t2 gnd 0.134f
C590 sensor_0.b.t10 gnd 0.127f
C591 sensor_0.b.t8 gnd 0.127f
C592 sensor_0.b.t16 gnd 0.0845f
C593 sensor_0.b.n11 gnd 0.0519f
C594 sensor_0.b.t3 gnd 0.00705f
C595 sensor_0.b.t11 gnd 0.00386f
C596 sensor_0.b.n12 gnd 0.138f
C597 sensor_0.b.t9 gnd 0.00386f
C598 sensor_0.b.n13 gnd 0.073f
C599 sensor_0.b.t17 gnd 0.00389f
C600 sensor_0.b.n14 gnd 0.0704f
C601 sensor_0.b.n15 gnd 0.0509f
C602 vd.t84 gnd 21.7f
C603 vd.t85 gnd 21.7f
C604 vd.t83 gnd 43.1f
C605 vd.n0 gnd 21.5f
C606 vd.n1 gnd 13.7f
C607 vd.t0 gnd 0.0573f
C608 vd.n2 gnd 17.5f
C609 vd.t55 gnd 0.00529f
C610 vd.t78 gnd 0.00264f
C611 vd.n3 gnd 0.00881f
C612 vd.t53 gnd 0.0301f
C613 vd.n4 gnd 0.191f
C614 vd.t66 gnd 0.00264f
C615 vd.t62 gnd 0.00264f
C616 vd.n5 gnd 0.0408f
C617 vd.n6 gnd 0.0645f
C618 vd.t58 gnd 0.00264f
C619 vd.t76 gnd 0.00264f
C620 vd.n7 gnd 0.0408f
C621 vd.n8 gnd 0.0539f
C622 vd.t74 gnd 0.00363f
C623 vd.n9 gnd 0.0826f
C624 vd.t64 gnd 0.00363f
C625 vd.n10 gnd 0.0782f
C626 vd.t60 gnd 0.00264f
C627 vd.t70 gnd 0.00264f
C628 vd.n11 gnd 0.0408f
C629 vd.n12 gnd 0.0488f
C630 vd.t68 gnd 0.00264f
C631 vd.t72 gnd 0.00264f
C632 vd.n13 gnd 0.0408f
C633 vd.n14 gnd 0.0445f
C634 vd.t12 gnd 0.00363f
C635 vd.n15 gnd 0.0869f
C636 vd.t10 gnd 0.00264f
C637 vd.t8 gnd 0.00264f
C638 vd.n16 gnd 0.0438f
C639 vd.n17 gnd 0.0486f
C640 vd.t6 gnd 0.00264f
C641 vd.t18 gnd 0.00264f
C642 vd.n18 gnd 0.0408f
C643 vd.n19 gnd 0.0539f
C644 vd.t16 gnd 0.00367f
C645 vd.n20 gnd 0.0913f
C646 vd.t14 gnd 0.00264f
C647 vd.t22 gnd 0.00264f
C648 vd.n21 gnd 0.0408f
C649 vd.n22 gnd 0.0437f
C650 vd.t4 gnd 0.00264f
C651 vd.t20 gnd 0.00264f
C652 vd.n23 gnd 0.0408f
C653 vd.n24 gnd 0.0368f
C654 vd.t48 gnd 0.00265f
C655 vd.t45 gnd 0.0301f
C656 vd.t2 gnd 0.00264f
C657 vd.t47 gnd 0.00264f
C658 vd.n25 gnd 0.00698f
C659 vd.n26 gnd 0.184f
C660 vd.t61 gnd 0.161f
C661 vd.t65 gnd 0.161f
C662 vd.t77 gnd 0.161f
C663 vd.t54 gnd 0.161f
C664 vd.n27 gnd 0.227f
C665 vd.n28 gnd 0.113f
C666 vd.t57 gnd 0.161f
C667 vd.t75 gnd 0.199f
C668 vd.t73 gnd 0.24f
C669 vd.t63 gnd 0.202f
C670 vd.t59 gnd 0.161f
C671 vd.t69 gnd 0.161f
C672 vd.t67 gnd 0.113f
C673 vd.n29 gnd 0.0806f
C674 vd.n30 gnd 0.0589f
C675 vd.n31 gnd 0.0589f
C676 vd.t71 gnd 0.106f
C677 vd.n32 gnd 0.118f
C678 vd.n33 gnd 0.118f
C679 vd.t5 gnd 0.161f
C680 vd.t7 gnd 0.161f
C681 vd.t9 gnd 0.161f
C682 vd.t11 gnd 0.144f
C683 vd.n34 gnd 0.121f
C684 vd.n35 gnd 0.0497f
C685 vd.n36 gnd 0.0493f
C686 vd.t17 gnd 0.199f
C687 vd.t15 gnd 0.234f
C688 vd.t13 gnd 0.196f
C689 vd.t21 gnd 0.161f
C690 vd.t3 gnd 0.161f
C691 vd.t19 gnd 0.115f
C692 vd.t1 gnd 0.106f
C693 vd.n37 gnd 0.0806f
C694 vd.n38 gnd 0.0497f
C695 vd.n39 gnd 0.181f
C696 vd.n40 gnd 0.0688f
C697 vd.t46 gnd 0.1f
C698 vd.n41 gnd 0.0806f
C699 vd.n42 gnd 0.0147f
C700 vd.n43 gnd 0.0144f
C701 vd.n44 gnd 0.0532f
C702 vd.n45 gnd 0.0143f
C703 vd.n46 gnd 0.102f
C704 vd.n47 gnd 0.0142f
C705 vd.n48 gnd 0.00352f
C706 vd.n49 gnd 0.0108f
C707 vd.n50 gnd 6.74e-19
C708 vd.t33 gnd 0.00793f
C709 vd.n51 gnd 0.00188f
C710 vd.n52 gnd 0.0124f
C711 vd.n53 gnd 0.00255f
C712 vd.n54 gnd 0.0143f
C713 vd.n55 gnd 7.28e-19
C714 vd.n56 gnd 0.00522f
C715 vd.n57 gnd 0.0143f
C716 vd.t32 gnd 0.149f
C717 vd.n59 gnd 0.0142f
C718 vd.n60 gnd 0.00522f
C719 vd.n62 gnd 0.144f
C720 vd.n63 gnd 0.0191f
C721 vd.n64 gnd 0.0142f
C722 vd.n65 gnd 0.00581f
C723 vd.n66 gnd 0.0096f
C724 vd.n67 gnd 0.125f
C725 vd.n68 gnd 0.0097f
C726 vd.n69 gnd 0.00593f
C727 vd.n70 gnd 0.0151f
C728 vd.n71 gnd 0.0302f
C729 vd.n72 gnd 0.0153f
C730 vd.n73 gnd 0.00837f
C731 vd.n74 gnd 0.0461f
C732 vd.n75 gnd 0.00327f
C733 vd.n76 gnd 0.00883f
C734 vd.n77 gnd 0.00182f
C735 vd.n78 gnd 0.00237f
C736 vd.n79 gnd 0.00219f
C737 vd.n80 gnd 0.0106f
C738 vd.n81 gnd 0.014f
C739 vd.n82 gnd 0.135f
C740 vd.t51 gnd 0.00556f
C741 vd.t52 gnd 0.00552f
C742 vd.t25 gnd 0.0058f
C743 vd.n83 gnd 0.0893f
C744 vd.t49 gnd 0.0924f
C745 vd.n84 gnd 0.0732f
C746 vd.n85 gnd 0.109f
C747 vd.n86 gnd 0.0576f
C748 vd.n87 gnd 0.291f
C749 vd.n88 gnd 0.232f
C750 vd.n89 gnd 0.019f
C751 vd.n90 gnd 0.019f
C752 vd.t80 gnd 0.0941f
C753 vd.t50 gnd 0.102f
C754 vd.t82 gnd 0.349f
C755 vd.n91 gnd 0.278f
C756 vd.n92 gnd 0.0108f
C757 vd.t36 gnd 0.156f
C758 vd.n93 gnd 0.196f
C759 vd.n94 gnd 0.0142f
C760 vd.n95 gnd 0.014f
C761 vd.n96 gnd 0.0119f
C762 vd.t44 gnd 0.00558f
C763 vd.t41 gnd 0.0924f
C764 vd.t43 gnd 0.00563f
C765 vd.t28 gnd 0.00588f
C766 vd.n97 gnd 0.102f
C767 vd.n98 gnd 0.0671f
C768 vd.n99 gnd 0.0801f
C769 vd.n100 gnd 0.00177f
C770 vd.t40 gnd 0.00529f
C771 vd.n101 gnd 0.0307f
C772 vd.t39 gnd 0.00556f
C773 vd.t31 gnd 0.00528f
C774 vd.t35 gnd 0.00528f
C775 vd.n102 gnd 0.0419f
C776 vd.n103 gnd 0.0544f
C777 vd.t37 gnd 0.0924f
C778 vd.n104 gnd 0.0612f
C779 vd.n105 gnd 0.00621f
C780 vd.n106 gnd 0.00285f
C781 vd.n107 gnd 0.051f
C782 vd.n108 gnd 0.0593f
C783 vd.n109 gnd 0.348f
C784 vd.t38 gnd 0.236f
C785 vd.n110 gnd 0.288f
C786 vd.n111 gnd 0.0224f
C787 vd.n112 gnd 0.0223f
C788 vd.t30 gnd 0.425f
C789 vd.t34 gnd 0.265f
C790 vd.n113 gnd 0.196f
C791 vd.n114 gnd 0.0141f
C792 vd.n115 gnd 0.0152f
C793 vd.n116 gnd 0.119f
C794 vd.n117 gnd 0.142f
C795 vd.t29 gnd 0.103f
C796 vd.t27 gnd 0.0819f
C797 vd.n118 gnd 0.0846f
C798 vd.n119 gnd 0.0846f
C799 vd.n120 gnd 0.17f
C800 vd.n121 gnd 0.00604f
C801 vd.n122 gnd 0.00602f
C802 vd.t81 gnd 0.252f
C803 vd.n123 gnd 0.29f
C804 vd.n124 gnd 0.0173f
C805 vd.n125 gnd 0.0171f
C806 vd.t56 gnd 0.137f
C807 vd.t26 gnd 0.273f
C808 vd.t42 gnd 0.173f
C809 vd.n126 gnd 0.118f
C810 vd.n127 gnd 0.0115f
C811 vd.n128 gnd 0.0125f
C812 vd.n129 gnd 0.117f
C813 vd.n130 gnd 0.293f
C814 vd.n131 gnd 0.00929f
C815 vd.n132 gnd 0.00918f
C816 vd.t24 gnd 0.196f
C817 vd.t23 gnd 0.193f
C818 vd.t79 gnd 0.296f
C819 vd.n133 gnd 0.196f
C820 vd.n134 gnd 0.0132f
C821 vd.n135 gnd 0.0143f
C822 vd.n136 gnd 0.166f
C823 vd.n137 gnd 0.0961f
C824 vd.n138 gnd 0.563f
C825 vd.n139 gnd 1.81f
C826 vd.n140 gnd 5.37f
C827 vd.n141 gnd 4.9f
C828 vd.n142 gnd 0.461f
C829 buffer_0.a.n0 gnd 1.52f
C830 buffer_0.a.n1 gnd 1.5f
C831 buffer_0.a.t6 gnd 0.0207f
C832 buffer_0.a.t21 gnd 0.514f
C833 buffer_0.a.t22 gnd 0.509f
C834 buffer_0.a.n2 gnd 0.575f
C835 buffer_0.a.t23 gnd 0.509f
C836 buffer_0.a.n3 gnd 0.295f
C837 buffer_0.a.t24 gnd 0.509f
C838 buffer_0.a.n4 gnd 0.295f
C839 buffer_0.a.t19 gnd 0.509f
C840 buffer_0.a.n5 gnd 0.295f
C841 buffer_0.a.t5 gnd 0.509f
C842 buffer_0.a.t20 gnd 0.509f
C843 buffer_0.a.t17 gnd 0.509f
C844 buffer_0.a.t25 gnd 0.509f
C845 buffer_0.a.t18 gnd 0.509f
C846 buffer_0.a.t26 gnd 0.514f
C847 buffer_0.a.n6 gnd 0.574f
C848 buffer_0.a.n7 gnd 0.295f
C849 buffer_0.a.n8 gnd 0.295f
C850 buffer_0.a.n9 gnd 0.311f
C851 buffer_0.a.n10 gnd 0.291f
C852 buffer_0.a.n11 gnd 0.0789f
C853 buffer_0.a.n12 gnd 0.352f
C854 buffer_0.a.t0 gnd 0.393f
C855 buffer_0.a.t1 gnd 0.0421f
C856 buffer_0.a.t13 gnd 0.0207f
C857 buffer_0.a.t15 gnd 0.0207f
C858 buffer_0.a.t12 gnd 0.0207f
C859 buffer_0.a.n13 gnd 0.304f
C860 buffer_0.a.n14 gnd 0.582f
C861 buffer_0.a.t11 gnd 0.0207f
C862 buffer_0.a.t10 gnd 0.0207f
C863 buffer_0.a.n15 gnd 0.302f
C864 buffer_0.a.n16 gnd 0.515f
C865 buffer_0.a.t16 gnd 0.0207f
C866 buffer_0.a.t14 gnd 0.0207f
C867 buffer_0.a.n17 gnd 0.304f
C868 buffer_0.a.n18 gnd 0.384f
C869 buffer_0.a.t7 gnd 0.0207f
C870 buffer_0.a.t8 gnd 0.0207f
C871 buffer_0.a.n19 gnd 0.301f
C872 buffer_0.a.t2 gnd 0.398f
C873 buffer_0.a.t9 gnd 0.0207f
C874 buffer_0.a.t3 gnd 0.0207f
C875 buffer_0.a.t4 gnd 0.0207f
C876 buffer_0.a.n20 gnd 0.486f
C877 buffer_0.a.n21 gnd 0.293f
C878 out_buff.t0 gnd 0.0837f
C879 out_buff.t6 gnd 0.004f
C880 out_buff.t3 gnd 0.004f
C881 out_buff.n0 gnd 0.0547f
C882 out_buff.t20 gnd 0.004f
C883 out_buff.t15 gnd 0.004f
C884 out_buff.n1 gnd 0.0902f
C885 out_buff.t13 gnd 0.004f
C886 out_buff.t11 gnd 0.004f
C887 out_buff.n2 gnd 0.0619f
C888 out_buff.n3 gnd 0.0803f
C889 out_buff.t19 gnd 0.0055f
C890 out_buff.n4 gnd 0.124f
C891 out_buff.t14 gnd 0.004f
C892 out_buff.t12 gnd 0.004f
C893 out_buff.n5 gnd 0.0619f
C894 out_buff.t17 gnd 0.004f
C895 out_buff.t16 gnd 0.004f
C896 out_buff.n6 gnd 0.0664f
C897 out_buff.t18 gnd 0.00938f
C898 out_buff.n7 gnd 0.172f
C899 out_buff.n8 gnd 0.0558f
C900 out_buff.n9 gnd 0.083f
C901 out_buff.t2 gnd 0.004f
C902 out_buff.t4 gnd 0.004f
C903 out_buff.n10 gnd 0.0592f
C904 out_buff.t9 gnd 0.004f
C905 out_buff.t10 gnd 0.004f
C906 out_buff.n11 gnd 0.0547f
C907 out_buff.t1 gnd 0.004f
C908 out_buff.t5 gnd 0.004f
C909 out_buff.n12 gnd 0.0539f
C910 out_buff.t7 gnd 0.004f
C911 out_buff.t8 gnd 0.004f
C912 out_buff.n13 gnd 0.103f
C913 out_buff.n14 gnd 0.114f
C914 out_buff.n15 gnd 0.1f
C915 out_buff.n16 gnd 0.0645f
C916 out_buff.n17 gnd 0.0952f
C917 out_buff.n18 gnd 0.0571f
C918 out_buff.t28 gnd 49.8f
C919 out_buff.n19 gnd 0.209f
C920 out_buff.t25 gnd 0.0757f
C921 out_buff.t24 gnd 0.0823f
C922 out_buff.t23 gnd 0.0761f
C923 out_buff.n20 gnd 0.149f
C924 out_buff.t30 gnd 0.0774f
C925 out_buff.n21 gnd 0.0768f
C926 out_buff.t29 gnd 0.0766f
C927 out_buff.n22 gnd 0.078f
C928 out_buff.t21 gnd 0.0764f
C929 out_buff.n23 gnd 0.0775f
C930 out_buff.t26 gnd 0.0751f
C931 out_buff.n24 gnd 0.0805f
C932 out_buff.t27 gnd 0.0756f
C933 out_buff.n25 gnd 0.0797f
C934 out_buff.t31 gnd 0.0771f
C935 out_buff.n26 gnd 0.0776f
C936 out_buff.t22 gnd 0.0769f
C937 out_buff.n27 gnd 0.0774f
C938 out_buff.n28 gnd 0.116f
C939 out_buff.n29 gnd 0.14f
C940 out_buff.n30 gnd 0.392f
*.ends




**** end user architecture code
x1 vd out l0
.ends


* expanding   symbol:  /foss/designs/temp-sensor/ask_modulator/xschem/l0.sym # of pins=2
** sym_path: /foss/designs/temp-sensor/ask_modulator/xschem/l0.sym
** sch_path: /foss/designs/temp-sensor/ask_modulator/xschem/l0.sch
.subckt l0 p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 993p m=1
Cs1 p1 net1 58.53f m=1
Cs2 p2 net2 52.93f m=1
Rs1 net1 GND 24.1 m=1
Rs2 net2 GND 22.94 m=1
R1 p2 net3 3.443 m=1
.ends

.GLOBAL GND
.end
