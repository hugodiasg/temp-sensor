magic
tech sky130A
magscale 1 2
timestamp 1655684427
<< nwell >>
rect -554 -1019 554 1019
<< pmos >>
rect -358 -800 -158 800
rect -100 -800 100 800
rect 158 -800 358 800
<< pdiff >>
rect -416 788 -358 800
rect -416 -788 -404 788
rect -370 -788 -358 788
rect -416 -800 -358 -788
rect -158 788 -100 800
rect -158 -788 -146 788
rect -112 -788 -100 788
rect -158 -800 -100 -788
rect 100 788 158 800
rect 100 -788 112 788
rect 146 -788 158 788
rect 100 -800 158 -788
rect 358 788 416 800
rect 358 -788 370 788
rect 404 -788 416 788
rect 358 -800 416 -788
<< pdiffc >>
rect -404 -788 -370 788
rect -146 -788 -112 788
rect 112 -788 146 788
rect 370 -788 404 788
<< nsubdiff >>
rect -518 949 -422 983
rect 422 949 518 983
rect -518 887 -484 949
rect 484 887 518 949
rect -518 -949 -484 -887
rect 484 -949 518 -887
rect -518 -983 -422 -949
rect 422 -983 518 -949
<< nsubdiffcont >>
rect -422 949 422 983
rect -518 -887 -484 887
rect 484 -887 518 887
rect -422 -983 422 -949
<< poly >>
rect -358 881 -158 897
rect -358 847 -342 881
rect -174 847 -158 881
rect -358 800 -158 847
rect -100 881 100 897
rect -100 847 -84 881
rect 84 847 100 881
rect -100 800 100 847
rect 158 881 358 897
rect 158 847 174 881
rect 342 847 358 881
rect 158 800 358 847
rect -358 -847 -158 -800
rect -358 -881 -342 -847
rect -174 -881 -158 -847
rect -358 -897 -158 -881
rect -100 -847 100 -800
rect -100 -881 -84 -847
rect 84 -881 100 -847
rect -100 -897 100 -881
rect 158 -847 358 -800
rect 158 -881 174 -847
rect 342 -881 358 -847
rect 158 -897 358 -881
<< polycont >>
rect -342 847 -174 881
rect -84 847 84 881
rect 174 847 342 881
rect -342 -881 -174 -847
rect -84 -881 84 -847
rect 174 -881 342 -847
<< locali >>
rect -518 949 -422 983
rect 422 949 518 983
rect -518 887 -484 949
rect 484 887 518 949
rect -358 847 -342 881
rect -174 847 -158 881
rect -100 847 -84 881
rect 84 847 100 881
rect 158 847 174 881
rect 342 847 358 881
rect -404 788 -370 804
rect -404 -804 -370 -788
rect -146 788 -112 804
rect -146 -804 -112 -788
rect 112 788 146 804
rect 112 -804 146 -788
rect 370 788 404 804
rect 370 -804 404 -788
rect -358 -881 -342 -847
rect -174 -881 -158 -847
rect -100 -881 -84 -847
rect 84 -881 100 -847
rect 158 -881 174 -847
rect 342 -881 358 -847
rect -518 -949 -484 -887
rect 484 -949 518 -887
rect -518 -983 -422 -949
rect 422 -983 518 -949
<< viali >>
rect -342 847 -174 881
rect -84 847 84 881
rect 174 847 342 881
rect -404 141 -370 771
rect -146 -315 -112 315
rect 112 141 146 771
rect 370 -315 404 315
rect -342 -881 -174 -847
rect -84 -881 84 -847
rect 174 -881 342 -847
<< metal1 >>
rect -354 881 -162 887
rect -354 847 -342 881
rect -174 847 -162 881
rect -354 841 -162 847
rect -96 881 96 887
rect -96 847 -84 881
rect 84 847 96 881
rect -96 841 96 847
rect 162 881 354 887
rect 162 847 174 881
rect 342 847 354 881
rect 162 841 354 847
rect -410 771 -364 783
rect -410 141 -404 771
rect -370 141 -364 771
rect 106 771 152 783
rect -410 129 -364 141
rect -152 315 -106 327
rect -152 -315 -146 315
rect -112 -315 -106 315
rect 106 141 112 771
rect 146 141 152 771
rect 106 129 152 141
rect 364 315 410 327
rect -152 -327 -106 -315
rect 364 -315 370 315
rect 404 -315 410 315
rect 364 -327 410 -315
rect -354 -847 -162 -841
rect -354 -881 -342 -847
rect -174 -881 -162 -847
rect -354 -887 -162 -881
rect -96 -847 96 -841
rect -96 -881 -84 -847
rect 84 -881 96 -847
rect -96 -887 96 -881
rect 162 -847 354 -841
rect 162 -881 174 -847
rect 342 -881 354 -847
rect 162 -887 354 -881
<< properties >>
string FIXED_BBOX -501 -966 501 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
