magic
tech sky130A
magscale 1 2
timestamp 1644351742
<< metal4 >>
rect -2549 7469 2549 7510
rect -2549 2611 2293 7469
rect 2529 2611 2549 7469
rect -2549 2570 2549 2611
rect -2549 2429 2549 2470
rect -2549 -2429 2293 2429
rect 2529 -2429 2549 2429
rect -2549 -2470 2549 -2429
rect -2549 -2611 2549 -2570
rect -2549 -7469 2293 -2611
rect 2529 -7469 2549 -2611
rect -2549 -7510 2549 -7469
<< via4 >>
rect 2293 2611 2529 7469
rect 2293 -2429 2529 2429
rect 2293 -7469 2529 -2611
<< mimcap2 >>
rect -2449 7370 2291 7410
rect -2449 2710 -2059 7370
rect 1901 2710 2291 7370
rect -2449 2670 2291 2710
rect -2449 2330 2291 2370
rect -2449 -2330 -2059 2330
rect 1901 -2330 2291 2330
rect -2449 -2370 2291 -2330
rect -2449 -2710 2291 -2670
rect -2449 -7370 -2059 -2710
rect 1901 -7370 2291 -2710
rect -2449 -7410 2291 -7370
<< mimcap2contact >>
rect -2059 2710 1901 7370
rect -2059 -2330 1901 2330
rect -2059 -7370 1901 -2710
<< metal5 >>
rect -239 7394 81 7560
rect 2251 7469 2571 7560
rect -2083 7370 1925 7394
rect -2083 2710 -2059 7370
rect 1901 2710 1925 7370
rect -2083 2686 1925 2710
rect -239 2354 81 2686
rect 2251 2611 2293 7469
rect 2529 2611 2571 7469
rect 2251 2429 2571 2611
rect -2083 2330 1925 2354
rect -2083 -2330 -2059 2330
rect 1901 -2330 1925 2330
rect -2083 -2354 1925 -2330
rect -239 -2686 81 -2354
rect 2251 -2429 2293 2429
rect 2529 -2429 2571 2429
rect 2251 -2611 2571 -2429
rect -2083 -2710 1925 -2686
rect -2083 -7370 -2059 -2710
rect 1901 -7370 1925 -2710
rect -2083 -7394 1925 -7370
rect -239 -7560 81 -7394
rect 2251 -7469 2293 -2611
rect 2529 -7469 2571 -2611
rect 2251 -7560 2571 -7469
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2549 2570 2391 7510
string parameters w 23.7 l 23.7 val 1.141k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 85
string library sky130
<< end >>
