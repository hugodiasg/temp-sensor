magic
tech sky130A
magscale 1 2
timestamp 1645798939
<< metal4 >>
rect -2829 11109 2829 11150
rect -2829 5691 2573 11109
rect 2809 5691 2829 11109
rect -2829 5650 2829 5691
rect -2829 5509 2829 5550
rect -2829 91 2573 5509
rect 2809 91 2829 5509
rect -2829 50 2829 91
rect -2829 -91 2829 -50
rect -2829 -5509 2573 -91
rect 2809 -5509 2829 -91
rect -2829 -5550 2829 -5509
rect -2829 -5691 2829 -5650
rect -2829 -11109 2573 -5691
rect 2809 -11109 2829 -5691
rect -2829 -11150 2829 -11109
<< via4 >>
rect 2573 5691 2809 11109
rect 2573 91 2809 5509
rect 2573 -5509 2809 -91
rect 2573 -11109 2809 -5691
<< mimcap2 >>
rect -2729 11010 2571 11050
rect -2729 5790 -2167 11010
rect 2009 5790 2571 11010
rect -2729 5750 2571 5790
rect -2729 5410 2571 5450
rect -2729 190 -2167 5410
rect 2009 190 2571 5410
rect -2729 150 2571 190
rect -2729 -190 2571 -150
rect -2729 -5410 -2167 -190
rect 2009 -5410 2571 -190
rect -2729 -5450 2571 -5410
rect -2729 -5790 2571 -5750
rect -2729 -11010 -2167 -5790
rect 2009 -11010 2571 -5790
rect -2729 -11050 2571 -11010
<< mimcap2contact >>
rect -2167 5790 2009 11010
rect -2167 190 2009 5410
rect -2167 -5410 2009 -190
rect -2167 -11010 2009 -5790
<< metal5 >>
rect -239 11034 81 11200
rect 2531 11109 2851 11200
rect -2191 11010 2033 11034
rect -2191 5790 -2167 11010
rect 2009 5790 2033 11010
rect -2191 5766 2033 5790
rect -239 5434 81 5766
rect 2531 5691 2573 11109
rect 2809 5691 2851 11109
rect 2531 5509 2851 5691
rect -2191 5410 2033 5434
rect -2191 190 -2167 5410
rect 2009 190 2033 5410
rect -2191 166 2033 190
rect -239 -166 81 166
rect 2531 91 2573 5509
rect 2809 91 2851 5509
rect 2531 -91 2851 91
rect -2191 -190 2033 -166
rect -2191 -5410 -2167 -190
rect 2009 -5410 2033 -190
rect -2191 -5434 2033 -5410
rect -239 -5766 81 -5434
rect 2531 -5509 2573 -91
rect 2809 -5509 2851 -91
rect 2531 -5691 2851 -5509
rect -2191 -5790 2033 -5766
rect -2191 -11010 -2167 -5790
rect 2009 -11010 2033 -5790
rect -2191 -11034 2033 -11010
rect -239 -11200 81 -11034
rect 2531 -11109 2573 -5691
rect 2809 -11109 2851 -5691
rect 2531 -11200 2851 -11109
<< properties >>
string FIXED_BBOX -2829 5650 2671 11150
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 26.5 l 26.5 val 1.424k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
