magic
tech sky130A
magscale 1 2
timestamp 1643598004
<< metal3 >>
rect -2121 2043 2120 2071
rect -2121 -2043 2036 2043
rect 2100 -2043 2120 2043
rect -2121 -2071 2120 -2043
<< via3 >>
rect 2036 -2043 2100 2043
<< mimcap >>
rect -2021 1931 1921 1971
rect -2021 -1931 -1981 1931
rect 1881 -1931 1921 1931
rect -2021 -1971 1921 -1931
<< mimcapcontact >>
rect -1981 -1931 1881 1931
<< metal4 >>
rect 2020 2043 2116 2059
rect -1982 1931 1882 1932
rect -1982 -1931 -1981 1931
rect 1881 -1931 1882 1931
rect -1982 -1932 1882 -1931
rect 2020 -2043 2036 2043
rect 2100 -2043 2116 2043
rect 2020 -2059 2116 -2043
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -2121 -2071 2021 2071
string parameters w 19.713 l 19.713 val 792.186 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
