magic
tech sky130A
magscale 1 2
timestamp 1644598236
use 1  1_0
timestamp 1644598236
transform 1 0 -116 0 1 -141
box 0 0 16000 16800
<< labels >>
flabel space 5963 16400 5963 16400 0 FreeSans 1600 0 0 0 p2
port 1 nsew
flabel space 335 15618 335 15618 0 FreeSans 1600 0 0 0 p1
port 0 nsew
<< end >>
