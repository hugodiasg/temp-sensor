magic
tech sky130A
magscale 1 2
timestamp 1646064585
<< metal4 >>
rect -2770 8132 2770 8173
rect -2770 2832 2514 8132
rect 2750 2832 2770 8132
rect -2770 2791 2770 2832
rect -2770 2650 2770 2691
rect -2770 -2650 2514 2650
rect 2750 -2650 2770 2650
rect -2770 -2691 2770 -2650
rect -2770 -2832 2770 -2791
rect -2770 -8132 2514 -2832
rect 2750 -8132 2770 -2832
rect -2770 -8173 2770 -8132
<< via4 >>
rect 2514 2832 2750 8132
rect 2514 -2650 2750 2650
rect 2514 -8132 2750 -2832
<< mimcap2 >>
rect -2670 8033 2512 8073
rect -2670 2931 -2120 8033
rect 1962 2931 2512 8033
rect -2670 2891 2512 2931
rect -2670 2551 2512 2591
rect -2670 -2551 -2120 2551
rect 1962 -2551 2512 2551
rect -2670 -2591 2512 -2551
rect -2670 -2931 2512 -2891
rect -2670 -8033 -2120 -2931
rect 1962 -8033 2512 -2931
rect -2670 -8073 2512 -8033
<< mimcap2contact >>
rect -2120 2931 1962 8033
rect -2120 -2551 1962 2551
rect -2120 -8033 1962 -2931
<< metal5 >>
rect -239 8057 81 8223
rect 2472 8132 2792 8223
rect -2144 8033 1986 8057
rect -2144 2931 -2120 8033
rect 1962 2931 1986 8033
rect -2144 2907 1986 2931
rect -239 2575 81 2907
rect 2472 2832 2514 8132
rect 2750 2832 2792 8132
rect 2472 2650 2792 2832
rect -2144 2551 1986 2575
rect -2144 -2551 -2120 2551
rect 1962 -2551 1986 2551
rect -2144 -2575 1986 -2551
rect -239 -2907 81 -2575
rect 2472 -2650 2514 2650
rect 2750 -2650 2792 2650
rect 2472 -2832 2792 -2650
rect -2144 -2931 1986 -2907
rect -2144 -8033 -2120 -2931
rect 1962 -8033 1986 -2931
rect -2144 -8057 1986 -8033
rect -239 -8223 81 -8057
rect 2472 -8132 2514 -2832
rect 2750 -8132 2792 -2832
rect 2472 -8223 2792 -8132
<< properties >>
string FIXED_BBOX -2770 2791 2612 8173
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.911 l 25.911 val 1.362k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
