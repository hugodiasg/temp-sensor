* NGSPICE file created from sigma-delta.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_EFDHR4 a_n33_n397# a_n73_n300# a_15_n300# w_n211_n519#
X0 a_15_n300# a_n33_n397# a_n73_n300# w_n211_n519# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VPWR Q Q_N VNB VPB
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=1.5393e+12p ps=1.452e+07u w=1e+06u l=150000u
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.2225e+12p pd=1.139e+07u as=0p ps=0u w=420000u l=150000u
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_EK42PW a_380_n1032# a_48_600# a_380_600# a_n450_n1032#
+ a_214_n1032# a_214_600# a_48_n1032# a_n284_600# a_n118_600# a_n580_n1162# a_n284_n1032#
+ a_n450_600# a_n118_n1032#
X0 a_380_n1032# a_380_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X1 a_214_n1032# a_214_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X2 a_n284_n1032# a_n284_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X3 a_n450_n1032# a_n450_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X4 a_48_n1032# a_48_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X5 a_n118_n1032# a_n118_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_X78HBF a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_A4KLY5 c1_n2770_n2720# m3_n2870_n2820#
X0 c1_n2770_n2720# m3_n2870_n2820# sky130_fd_pr__cap_mim_m3_1 l=2.72e+07u w=2.72e+07u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_ARMGAU a_380_n1032# a_48_600# a_380_600# a_n450_n1032#
+ a_214_n1032# a_214_600# a_48_n1032# a_n284_600# a_n118_600# a_n580_n1162# a_n284_n1032#
+ a_n450_600# a_n118_n1032#
X0 a_380_n1032# a_380_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X1 a_214_n1032# a_214_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X2 a_n284_n1032# a_n284_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X3 a_n450_n1032# a_n450_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X4 a_48_n1032# a_48_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X5 a_n118_n1032# a_n118_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
.ends

.subckt sigma-delta in vpwr out clk reset_b_dff gnd vd
Xsky130_fd_pr__pfet_01v8_EFDHR4_0 in_comp vd out_comp vd sky130_fd_pr__pfet_01v8_EFDHR4
Xx1 clk out_comp reset_b_dff gnd vpwr Q out gnd vpwr sky130_fd_sc_hd__dfrbp_1
XXR2 Q m1_n1710_5800# m1_n1400_5790# in_comp m1_n1550_4170# m1_n1400_5790# m1_n1550_4170#
+ m1_n2050_5780# m1_n1710_5800# gnd m1_n1890_4160# m1_n2050_5780# m1_n1890_4160# sky130_fd_pr__res_xhigh_po_0p35_EK42PW
XXN1 gnd in_comp out_comp gnd sky130_fd_pr__nfet_01v8_X78HBF
XXC1 in_comp gnd sky130_fd_pr__cap_mim_m3_1_A4KLY5
Xsky130_fd_pr__res_xhigh_po_0p35_ARMGAU_0 in_comp m1_n3250_5800# m1_n2930_5790# in
+ m1_n3070_4170# m1_n2930_5790# m1_n3070_4170# m1_n3590_5800# m1_n3250_5800# gnd m1_n3420_4160#
+ m1_n3590_5800# m1_n3420_4160# sky130_fd_pr__res_xhigh_po_0p35_ARMGAU
.ends

