magic
tech sky130A
magscale 1 2
timestamp 1645495691
<< metal4 >>
rect 32200 68519 33478 71480
rect 32199 67241 33478 68519
rect 32200 67240 33478 67241
<< metal5 >>
rect 32200 68918 70200 70200
rect 32200 68519 33478 68520
rect 32199 67241 33478 68519
rect 32200 33478 33478 67241
rect 68918 33478 70200 68918
rect 32200 32200 70200 33478
<< end >>
