magic
tech sky130A
magscale 1 2
timestamp 1645036902
<< metal4 >>
rect -2514 7364 2514 7405
rect -2514 2576 2258 7364
rect 2494 2576 2514 7364
rect -2514 2535 2514 2576
rect -2514 2394 2514 2435
rect -2514 -2394 2258 2394
rect 2494 -2394 2514 2394
rect -2514 -2435 2514 -2394
rect -2514 -2576 2514 -2535
rect -2514 -7364 2258 -2576
rect 2494 -7364 2514 -2576
rect -2514 -7405 2514 -7364
<< via4 >>
rect 2258 2576 2494 7364
rect 2258 -2394 2494 2394
rect 2258 -7364 2494 -2576
<< mimcap2 >>
rect -2414 7265 2256 7305
rect -2414 2675 -1915 7265
rect 1757 2675 2256 7265
rect -2414 2635 2256 2675
rect -2414 2295 2256 2335
rect -2414 -2295 -1915 2295
rect 1757 -2295 2256 2295
rect -2414 -2335 2256 -2295
rect -2414 -2675 2256 -2635
rect -2414 -7265 -1915 -2675
rect 1757 -7265 2256 -2675
rect -2414 -7305 2256 -7265
<< mimcap2contact >>
rect -1915 2675 1757 7265
rect -1915 -2295 1757 2295
rect -1915 -7265 1757 -2675
<< metal5 >>
rect -239 7289 81 7455
rect 2216 7364 2536 7455
rect -1939 7265 1781 7289
rect -1939 2675 -1915 7265
rect 1757 2675 1781 7265
rect -1939 2651 1781 2675
rect -239 2319 81 2651
rect 2216 2576 2258 7364
rect 2494 2576 2536 7364
rect 2216 2394 2536 2576
rect -1939 2295 1781 2319
rect -1939 -2295 -1915 2295
rect 1757 -2295 1781 2295
rect -1939 -2319 1781 -2295
rect -239 -2651 81 -2319
rect 2216 -2394 2258 2394
rect 2494 -2394 2536 2394
rect 2216 -2576 2536 -2394
rect -1939 -2675 1781 -2651
rect -1939 -7265 -1915 -2675
rect 1757 -7265 1781 -2675
rect -1939 -7289 1781 -7265
rect -239 -7455 81 -7289
rect 2216 -7364 2258 -2576
rect 2494 -7364 2536 -2576
rect 2216 -7455 2536 -7364
<< properties >>
string FIXED_BBOX -2514 2535 2356 7405
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.35 l 23.35 val 1.108k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
