magic
tech sky130A
magscale 1 2
timestamp 1644168429
<< metal1 >>
rect 15700 6500 16300 8700
rect 11800 6400 16300 6500
rect 11800 5600 11900 6400
rect 12700 5600 16300 6400
rect 11800 5400 16300 5600
rect 14980 1960 15380 5400
rect 15700 3400 16300 5400
rect 16600 6500 17200 8700
rect 16600 6400 20700 6500
rect 16600 5600 19800 6400
rect 20600 5600 20700 6400
rect 16600 5400 20700 5600
rect 16600 3400 17200 5400
rect 15780 2700 17480 3300
rect 16700 2400 17480 2700
rect 14980 1180 16320 1960
rect 16440 1800 17480 2400
rect 14980 -1120 15380 1180
rect 16200 -1120 16600 820
rect 17080 -1120 17480 1800
rect 18700 -1120 19100 5400
rect 15080 -1320 15280 -1120
rect 16300 -1320 16500 -1120
rect 17160 -1320 17360 -1120
rect 18800 -1320 19000 -1120
<< via1 >>
rect 11900 5600 12700 6400
rect 19800 5600 20600 6400
<< metal2 >>
rect 11800 6400 12800 6500
rect 11800 5600 11900 6400
rect 12700 5600 12800 6400
rect 11800 5400 12800 5600
rect 19700 6400 20700 6500
rect 19700 5600 19800 6400
rect 20600 5600 20700 6400
rect 19700 5400 20700 5600
<< via2 >>
rect 11900 5600 12700 6400
rect 19800 5600 20600 6400
<< metal3 >>
rect 11800 6400 12800 6500
rect 11800 5600 11900 6400
rect 12700 5600 12800 6400
rect 11800 5400 12800 5600
rect 19700 6400 20700 6500
rect 19700 5600 19800 6400
rect 20600 5600 20700 6400
rect 19700 5400 20700 5600
<< via3 >>
rect 11900 5600 12700 6400
rect 19800 5600 20600 6400
<< metal4 >>
rect 11800 27100 39100 28100
rect 11800 6400 12800 27100
rect 16200 24100 17100 27100
rect 38100 19100 39100 27100
rect 11800 5600 11900 6400
rect 12700 5600 12800 6400
rect 11800 5400 12800 5600
rect 19700 6400 20700 6500
rect 19700 5600 19800 6400
rect 20600 5600 20700 6400
rect 19700 5400 20700 5600
<< via4 >>
rect 30100 19200 30800 19980
rect 19800 5600 20600 6400
<< metal5 >>
rect 16200 25500 34900 26500
rect 16200 24100 17100 25500
rect 19700 6400 20700 25500
rect 30076 19980 30824 20004
rect 30076 19200 30100 19980
rect 30800 19200 30824 19980
rect 30076 19176 30824 19200
rect 19700 5600 19800 6400
rect 20600 5600 20700 6400
rect 19700 5400 20700 5600
use sky130_fd_pr__nfet_g5v0d10v5_FLFTBY  XM2
timestamp 1644164861
transform -1 0 16398 0 1 1688
box -278 -1128 278 1128
use sky130_fd_pr__res_high_po_5p73_CAGT5B  XR0
timestamp 1644161670
transform 0 1 16454 -1 0 6030
box -2830 -654 2830 654
use l0  l0_0
timestamp 1644072167
transform 1 0 21200 0 1 10300
box 0 0 17200 16200
use sky130_fd_pr__cap_mim_m3_2_U2MGMH  sky130_fd_pr__cap_mim_m3_2_U2MGMH_0
timestamp 1644161670
transform 1 0 16579 0 1 17150
box -2579 -7650 2601 7650
<< labels >>
flabel metal1 16300 -1320 16500 -1120 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 15080 -1320 15280 -1120 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 18800 -1320 19000 -1120 0 FreeSans 128 0 0 0 vd
port 3 nsew
flabel metal1 17160 -1320 17360 -1120 0 FreeSans 128 0 0 0 gnd
port 0 nsew
<< end >>
