magic
tech sky130A
magscale 1 2
timestamp 1656875210
<< pwell >>
rect -457 -708 457 708
<< mvnmos >>
rect -229 -450 -29 450
rect 29 -450 229 450
<< mvndiff >>
rect -287 438 -229 450
rect -287 -438 -275 438
rect -241 -438 -229 438
rect -287 -450 -229 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 229 438 287 450
rect 229 -438 241 438
rect 275 -438 287 438
rect 229 -450 287 -438
<< mvndiffc >>
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
<< mvpsubdiff >>
rect -421 660 421 672
rect -421 626 -313 660
rect 313 626 421 660
rect -421 614 421 626
rect -421 564 -363 614
rect -421 -564 -409 564
rect -375 -564 -363 564
rect 363 564 421 614
rect -421 -614 -363 -564
rect 363 -564 375 564
rect 409 -564 421 564
rect 363 -614 421 -564
rect -421 -626 421 -614
rect -421 -660 -313 -626
rect 313 -660 421 -626
rect -421 -672 421 -660
<< mvpsubdiffcont >>
rect -313 626 313 660
rect -409 -564 -375 564
rect 375 -564 409 564
rect -313 -660 313 -626
<< poly >>
rect -229 522 -29 538
rect -229 488 -213 522
rect -45 488 -29 522
rect -229 450 -29 488
rect 29 522 229 538
rect 29 488 45 522
rect 213 488 229 522
rect 29 450 229 488
rect -229 -488 -29 -450
rect -229 -522 -213 -488
rect -45 -522 -29 -488
rect -229 -538 -29 -522
rect 29 -488 229 -450
rect 29 -522 45 -488
rect 213 -522 229 -488
rect 29 -538 229 -522
<< polycont >>
rect -213 488 -45 522
rect 45 488 213 522
rect -213 -522 -45 -488
rect 45 -522 213 -488
<< locali >>
rect -409 626 -313 660
rect 313 626 409 660
rect -409 564 -375 626
rect 375 564 409 626
rect -229 488 -213 522
rect -45 488 -29 522
rect 29 488 45 522
rect 213 488 229 522
rect -275 438 -241 454
rect -275 -454 -241 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 241 438 275 454
rect 241 -454 275 -438
rect -229 -522 -213 -488
rect -45 -522 -29 -488
rect 29 -522 45 -488
rect 213 -522 229 -488
rect -409 -660 -375 -564
rect 375 -660 409 -564
<< viali >>
rect -213 488 -45 522
rect 45 488 213 522
rect -275 71 -241 421
rect -17 -175 17 175
rect 241 71 275 421
rect -213 -522 -45 -488
rect 45 -522 213 -488
rect -375 -660 -313 -626
rect -313 -660 313 -626
rect 313 -660 375 -626
<< metal1 >>
rect -225 522 -33 528
rect -225 488 -213 522
rect -45 488 -33 522
rect -225 482 -33 488
rect 33 522 225 528
rect 33 488 45 522
rect 213 488 225 522
rect 33 482 225 488
rect -281 421 -235 433
rect -281 71 -275 421
rect -241 71 -235 421
rect 235 421 281 433
rect -281 59 -235 71
rect -23 175 23 187
rect -23 -175 -17 175
rect 17 -175 23 175
rect 235 71 241 421
rect 275 71 281 421
rect 235 59 281 71
rect -23 -187 23 -175
rect -225 -488 -33 -482
rect -225 -522 -213 -488
rect -45 -522 -33 -488
rect -225 -528 -33 -522
rect 33 -488 225 -482
rect 33 -522 45 -488
rect 213 -522 225 -488
rect 33 -528 225 -522
rect -387 -626 387 -620
rect -387 -660 -375 -626
rect 375 -660 387 -626
rect -387 -666 387 -660
<< properties >>
string FIXED_BBOX -392 -643 392 643
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
