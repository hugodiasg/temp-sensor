magic
tech sky130A
magscale 1 2
timestamp 1656875000
<< nwell >>
rect -358 -897 358 897
<< mvpmos >>
rect -100 -600 100 600
<< mvpdiff >>
rect -158 588 -100 600
rect -158 -588 -146 588
rect -112 -588 -100 588
rect -158 -600 -100 -588
rect 100 588 158 600
rect 100 -588 112 588
rect 146 -588 158 588
rect 100 -600 158 -588
<< mvpdiffc >>
rect -146 -588 -112 588
rect 112 -588 146 588
<< mvnsubdiff >>
rect -292 819 292 831
rect -292 785 -184 819
rect 184 785 292 819
rect -292 773 292 785
rect -292 723 -234 773
rect -292 -723 -280 723
rect -246 -723 -234 723
rect 234 723 292 773
rect -292 -773 -234 -723
rect 234 -723 246 723
rect 280 -723 292 723
rect 234 -773 292 -723
rect -292 -785 292 -773
rect -292 -819 -184 -785
rect 184 -819 292 -785
rect -292 -831 292 -819
<< mvnsubdiffcont >>
rect -184 785 184 819
rect -280 -723 -246 723
rect 246 -723 280 723
rect -184 -819 184 -785
<< poly >>
rect -100 681 100 697
rect -100 647 -84 681
rect 84 647 100 681
rect -100 600 100 647
rect -100 -647 100 -600
rect -100 -681 -84 -647
rect 84 -681 100 -647
rect -100 -697 100 -681
<< polycont >>
rect -84 647 84 681
rect -84 -681 84 -647
<< locali >>
rect -280 785 -184 819
rect 184 785 280 819
rect -280 723 -246 785
rect 246 723 280 785
rect -100 647 -84 681
rect 84 647 100 681
rect -146 588 -112 604
rect -146 -604 -112 -588
rect 112 588 146 604
rect 112 -604 146 -588
rect -100 -681 -84 -647
rect 84 -681 100 -647
rect -280 -785 -246 -723
rect 246 -785 280 -723
rect -280 -819 -184 -785
rect 184 -819 280 -785
<< viali >>
rect -84 647 84 681
rect -146 -588 -112 588
rect 112 -588 146 588
rect -84 -681 84 -647
<< metal1 >>
rect -96 681 96 687
rect -96 647 -84 681
rect 84 647 96 681
rect -96 641 96 647
rect -152 588 -106 600
rect -152 -588 -146 588
rect -112 -588 -106 588
rect -152 -600 -106 -588
rect 106 588 152 600
rect 106 -588 112 588
rect 146 -588 152 588
rect 106 -600 152 -588
rect -96 -647 96 -641
rect -96 -681 -84 -647
rect 84 -681 96 -647
rect -96 -687 96 -681
<< properties >>
string FIXED_BBOX -263 -802 263 802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
