magic
tech sky130A
magscale 1 2
timestamp 1668740706
<< nwell >>
rect -296 -819 296 819
<< pmos >>
rect -100 -600 100 600
<< pdiff >>
rect -158 588 -100 600
rect -158 -588 -146 588
rect -112 -588 -100 588
rect -158 -600 -100 -588
rect 100 588 158 600
rect 100 -588 112 588
rect 146 -588 158 588
rect 100 -600 158 -588
<< pdiffc >>
rect -146 -588 -112 588
rect 112 -588 146 588
<< nsubdiff >>
rect -260 749 -164 783
rect 164 749 260 783
rect -260 687 -226 749
rect 226 687 260 749
rect -260 -749 -226 -687
rect 226 -749 260 -687
rect -260 -783 -164 -749
rect 164 -783 260 -749
<< nsubdiffcont >>
rect -164 749 164 783
rect -260 -687 -226 687
rect 226 -687 260 687
rect -164 -783 164 -749
<< poly >>
rect -100 681 100 697
rect -100 647 -84 681
rect 84 647 100 681
rect -100 600 100 647
rect -100 -647 100 -600
rect -100 -681 -84 -647
rect 84 -681 100 -647
rect -100 -697 100 -681
<< polycont >>
rect -84 647 84 681
rect -84 -681 84 -647
<< locali >>
rect -260 749 -164 783
rect 164 749 260 783
rect -260 687 -226 749
rect -100 647 -84 681
rect 84 647 100 681
rect -146 588 -112 604
rect -146 -604 -112 -588
rect 112 588 146 604
rect 112 -604 146 -588
rect -100 -681 -84 -647
rect 84 -681 100 -647
rect -260 -749 -226 -687
rect -260 -783 -164 -749
rect 164 -783 260 -749
<< viali >>
rect 226 687 260 749
rect -84 647 84 681
rect -146 -588 -112 588
rect 112 -588 146 588
rect -84 -681 84 -647
rect 226 -687 260 687
rect 226 -749 260 -687
<< metal1 >>
rect 220 749 266 761
rect -96 681 96 687
rect -96 647 -84 681
rect 84 647 96 681
rect -96 641 96 647
rect -152 588 -106 600
rect -152 -588 -146 588
rect -112 -588 -106 588
rect -152 -600 -106 -588
rect 106 588 152 600
rect 106 -588 112 588
rect 146 -588 152 588
rect 106 -600 152 -588
rect -96 -647 96 -641
rect -96 -681 -84 -647
rect 84 -681 96 -647
rect -96 -687 96 -681
rect 220 -749 226 749
rect 260 -749 266 749
rect 220 -761 266 -749
<< properties >>
string FIXED_BBOX -243 -766 243 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 100 viagl 0 viagt 0
<< end >>
