magic
tech sky130A
magscale 1 2
timestamp 1656876180
<< nwell >>
rect 460 9160 640 9380
<< metal1 >>
rect 2460 12760 2660 12960
rect 700 12700 4140 12760
rect 700 12020 760 12700
rect 1680 12020 1740 12700
rect 2320 12380 2380 12700
rect 2320 12320 3460 12380
rect 4080 12000 4140 12700
rect -100 11220 160 11420
rect 100 10860 160 11220
rect 980 11100 1100 11120
rect 980 11020 1000 11100
rect 1080 11080 1100 11100
rect 1080 11020 1420 11080
rect 2620 11040 2680 11420
rect 3140 11040 3200 11420
rect 3500 11040 3620 11060
rect 980 11000 1100 11020
rect 2620 10980 3520 11040
rect 3500 10960 3520 10980
rect 3600 10960 3620 11040
rect 400 10860 460 10960
rect 3500 10940 3620 10960
rect 100 10800 4380 10860
rect 4420 10520 4480 11000
rect -100 10460 100 10520
rect -100 10380 1640 10460
rect -100 10320 100 10380
rect 700 10040 760 10260
rect 980 10080 1100 10100
rect 1440 10080 1640 10380
rect 4420 10320 4840 10520
rect 980 10040 1000 10080
rect 680 10000 1000 10040
rect 1080 10040 1100 10080
rect 1080 10000 1420 10040
rect 680 9980 1420 10000
rect 4420 9940 4480 10320
rect 400 9540 520 9560
rect 400 9460 420 9540
rect 500 9460 520 9540
rect 400 9440 520 9460
rect 1000 9540 1120 9560
rect 1000 9460 1020 9540
rect 1100 9460 1120 9540
rect 2300 9540 3120 9600
rect 1000 9440 1120 9460
rect -100 9200 100 9280
rect 460 9200 640 9380
rect -100 9140 640 9200
rect -100 9080 100 9140
rect 1040 8920 1100 9440
rect 1680 9140 1740 9520
rect 2300 9140 2360 9540
rect 2660 9380 2860 9540
rect 2940 9380 3120 9540
rect 1680 9080 2360 9140
rect 2460 9260 4180 9320
rect 620 8860 1520 8920
rect -100 8360 100 8420
rect 540 8360 600 8820
rect 860 8600 920 8860
rect 1680 8820 1740 9080
rect 1240 8360 1300 8820
rect 1540 8740 1740 8820
rect 1540 8720 1760 8740
rect 1640 8640 1660 8720
rect 1740 8640 1760 8720
rect 1640 8620 1760 8640
rect 2460 8360 2520 9260
rect 3480 8840 3660 8860
rect 3480 8800 3500 8840
rect 2880 8740 3500 8800
rect 3480 8720 3500 8740
rect 3640 8760 3660 8840
rect 4180 8760 4380 8800
rect 3640 8720 4380 8760
rect 3480 8700 4380 8720
rect -100 8300 2520 8360
rect -100 8220 100 8300
rect 2460 8240 2580 8300
<< via1 >>
rect 1000 11020 1080 11100
rect 3520 10960 3600 11040
rect 1000 10000 1080 10080
rect 420 9460 500 9540
rect 1020 9460 1100 9540
rect 1660 8640 1740 8720
rect 3500 8720 3640 8840
<< metal2 >>
rect 980 11100 1100 11120
rect 980 11020 1000 11100
rect 1080 11020 1100 11100
rect 980 11000 1100 11020
rect 3500 11040 3620 11060
rect 1000 10100 1060 11000
rect 3500 10960 3520 11040
rect 3600 10960 3620 11040
rect 3500 10940 3620 10960
rect 980 10080 1100 10100
rect 980 10000 1000 10080
rect 1080 10000 1100 10080
rect 980 9980 1100 10000
rect 400 9540 520 9560
rect 400 9460 420 9540
rect 500 9520 520 9540
rect 1000 9540 1120 9560
rect 1000 9520 1020 9540
rect 500 9460 1020 9520
rect 1100 9460 1120 9540
rect 400 9440 520 9460
rect 1000 9440 1120 9460
rect 3520 8860 3580 10940
rect 3480 8840 3660 8860
rect 1640 8720 1760 8740
rect 1640 8640 1660 8720
rect 1740 8640 1760 8720
rect 3480 8720 3500 8840
rect 3640 8720 3660 8840
rect 3480 8700 3660 8720
rect 1640 8620 1760 8640
rect 1660 8140 1720 8620
rect 1600 8120 1800 8140
rect 1600 8020 1620 8120
rect 1780 8020 1800 8120
rect 1600 8000 1800 8020
<< via2 >>
rect 3500 8720 3640 8840
rect 1620 8020 1780 8120
<< metal3 >>
rect 3480 8840 3660 8860
rect 3480 8720 3500 8840
rect 3640 8720 3660 8840
rect 3480 8700 3660 8720
rect 1600 8120 1800 8140
rect 1600 8020 1620 8120
rect 1780 8020 1800 8120
rect 1600 7660 1800 8020
<< via3 >>
rect 3500 8720 3640 8840
<< metal4 >>
rect 3480 8840 3660 8860
rect 3480 8720 3500 8840
rect 3640 8720 3660 8840
rect 3480 7680 3660 8720
use sky130_fd_pr__cap_mim_m3_1_2NYK3R  XCC
timestamp 1656875000
transform 1 0 2450 0 1 5800
box -2250 -2200 2249 2200
use sky130_fd_pr__pfet_g5v0d10v5_GYM5UZ  XM1
timestamp 1656875158
transform 1 0 558 0 1 9737
box -358 -597 358 597
use sky130_fd_pr__pfet_g5v0d10v5_G8J5UZ  XM2
timestamp 1656875158
transform 1 0 1538 0 1 9737
box -358 -597 358 597
use sky130_fd_pr__nfet_g5v0d10v5_9YTB7P  XM3
timestamp 1656875158
transform 1 0 728 0 1 8718
box -328 -358 328 358
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  XM5
timestamp 1656875000
transform 1 0 558 0 1 11497
box -358 -897 358 897
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  XM6
timestamp 1656875000
transform 1 0 1538 0 1 11497
box -358 -897 358 897
use sky130_fd_pr__nfet_g5v0d10v5_G8BGHZ  XM7
timestamp 1656875210
transform 1 0 2897 0 1 8908
box -457 -708 457 708
use sky130_fd_pr__pfet_g5v0d10v5_8C84A7  XM8
timestamp 1656875000
transform 1 0 2905 0 1 11647
box -745 -1047 745 1047
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  XM10
timestamp 1656875000
transform 1 0 4278 0 1 11497
box -358 -897 358 897
use sky130_fd_pr__nfet_g5v0d10v5_9YTB7P  sky130_fd_pr__nfet_g5v0d10v5_9YTB7P_0
timestamp 1656875158
transform 1 0 1428 0 1 8718
box -328 -358 328 358
use sky130_fd_pr__pfet_g5v0d10v5_GYMD5T  sky130_fd_pr__pfet_g5v0d10v5_GYMD5T_0
timestamp 1656875000
transform 1 0 4278 0 1 9437
box -358 -897 358 897
<< labels >>
flabel metal1 2460 12760 2660 12960 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 -100 8220 100 8420 0 FreeSans 1600 0 0 0 vs
port 5 nsew
flabel metal1 4640 10320 4840 10520 0 FreeSans 1600 0 0 0 out
port 2 nsew
flabel metal1 -100 9080 100 9280 0 FreeSans 1600 0 0 0 in1
port 4 nsew
flabel metal1 -100 10320 100 10520 0 FreeSans 1600 0 0 0 in2
port 3 nsew
flabel metal1 -100 11220 100 11420 0 FreeSans 1600 0 0 0 ib
port 1 nsew
flabel space 1020 10580 1160 10620 0 FreeSans 800 0 0 0 b
flabel metal1 1080 9360 1080 9360 0 FreeSans 800 0 0 0 c
flabel metal2 1680 8220 1680 8220 0 FreeSans 800 0 0 0 d
flabel metal1 3400 8760 3400 8760 0 FreeSans 800 0 0 0 e
<< end >>
