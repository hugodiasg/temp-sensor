magic
tech sky130A
magscale 1 2
timestamp 1655684427
<< pwell >>
rect -2996 -310 2996 310
<< nmos >>
rect -2800 -100 2800 100
<< ndiff >>
rect -2858 88 -2800 100
rect -2858 -88 -2846 88
rect -2812 -88 -2800 88
rect -2858 -100 -2800 -88
rect 2800 88 2858 100
rect 2800 -88 2812 88
rect 2846 -88 2858 88
rect 2800 -100 2858 -88
<< ndiffc >>
rect -2846 -88 -2812 88
rect 2812 -88 2846 88
<< psubdiff >>
rect -2960 240 -2864 274
rect 2864 240 2960 274
rect -2960 178 -2926 240
rect 2926 178 2960 240
rect -2960 -240 -2926 -178
rect 2926 -240 2960 -178
rect -2960 -274 -2864 -240
rect 2864 -274 2960 -240
<< psubdiffcont >>
rect -2864 240 2864 274
rect -2960 -178 -2926 178
rect 2926 -178 2960 178
rect -2864 -274 2864 -240
<< poly >>
rect -2800 172 2800 188
rect -2800 138 -2784 172
rect 2784 138 2800 172
rect -2800 100 2800 138
rect -2800 -138 2800 -100
rect -2800 -172 -2784 -138
rect 2784 -172 2800 -138
rect -2800 -188 2800 -172
<< polycont >>
rect -2784 138 2784 172
rect -2784 -172 2784 -138
<< locali >>
rect -2960 240 -2864 274
rect 2864 240 2960 274
rect -2960 178 -2926 240
rect 2926 178 2960 240
rect -2800 138 -2784 172
rect 2784 138 2800 172
rect -2846 88 -2812 104
rect -2846 -104 -2812 -88
rect 2812 88 2846 104
rect 2812 -104 2846 -88
rect -2800 -172 -2784 -138
rect 2784 -172 2800 -138
rect -2960 -240 -2926 -178
rect 2926 -240 2960 -178
rect -2960 -274 -2864 -240
rect 2864 -274 2960 -240
<< viali >>
rect -2784 138 2784 172
rect -2846 1 -2812 71
rect 2812 -35 2846 35
rect -2784 -172 2784 -138
<< metal1 >>
rect -2796 172 2796 178
rect -2796 138 -2784 172
rect 2784 138 2796 172
rect -2796 132 2796 138
rect -2852 71 -2806 83
rect -2852 1 -2846 71
rect -2812 1 -2806 71
rect -2852 -11 -2806 1
rect 2806 35 2852 47
rect 2806 -35 2812 35
rect 2846 -35 2852 35
rect 2806 -47 2852 -35
rect -2796 -138 2796 -132
rect -2796 -172 -2784 -138
rect 2784 -172 2796 -138
rect -2796 -178 2796 -172
<< properties >>
string FIXED_BBOX -2943 -257 2943 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 28.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
