magic
tech sky130A
magscale 1 2
timestamp 1708093148
<< nwell >>
rect 207 3627 4233 5293
rect 5608 4802 11988 5542
rect 167 2307 3393 3373
rect 5635 2049 7001 4802
rect 10628 2042 11988 4802
rect 14320 1390 14740 1400
rect 14320 1160 16752 1390
rect 14560 1069 16752 1160
rect 17014 934 17436 1972
<< pwell >>
rect 0 160 3392 2080
rect 7308 4002 10500 4782
rect 7308 3562 8688 4002
rect 8708 3562 10500 4002
rect 7308 2582 10500 3562
rect 14360 2120 17552 5940
rect 15501 965 15687 1009
rect 16231 965 16702 1011
rect 14599 829 16702 965
rect 14627 791 14661 829
rect 17014 264 17436 884
<< nmos >>
rect 8690 4310 8720 4610
rect 8786 4310 8816 4610
rect 8882 4310 8912 4610
rect 8978 4310 9008 4610
rect 7666 3690 7866 3890
rect 7924 3690 8124 3890
rect 8182 3690 8382 3890
rect 8440 3690 8640 3890
rect 8826 2830 9026 3830
rect 9084 2830 9284 3830
rect 9342 2830 9542 3830
rect 9600 2830 9800 3830
rect 9858 2830 10058 3830
rect 10116 2830 10316 3830
rect 218 1672 418 1872
rect 598 1672 798 1872
rect 978 1672 1178 1872
rect 1358 1672 1558 1872
rect 1738 1672 1938 1872
rect 2118 1672 2318 1872
rect 2498 1672 2698 1872
rect 2878 1672 3078 1872
rect 218 1254 418 1454
rect 598 1254 798 1454
rect 978 1254 1178 1454
rect 1358 1254 1558 1454
rect 1738 1254 1938 1454
rect 2118 1254 2318 1454
rect 2498 1254 2698 1454
rect 2878 1254 3078 1454
rect 218 836 418 1036
rect 598 836 798 1036
rect 978 836 1178 1036
rect 1358 836 1558 1036
rect 1738 836 1938 1036
rect 2118 836 2318 1036
rect 2498 836 2698 1036
rect 2878 836 3078 1036
rect 218 418 418 618
rect 598 418 798 618
rect 978 418 1178 618
rect 1358 418 1558 618
rect 1738 418 1938 618
rect 2118 418 2318 618
rect 2498 418 2698 618
rect 2878 418 3078 618
rect 17210 474 17240 674
<< scnmos >>
rect 14677 855 14707 939
rect 14761 855 14791 939
rect 15016 855 15046 939
rect 15111 855 15141 927
rect 15207 855 15237 927
rect 15373 855 15403 939
rect 15445 855 15475 939
rect 15577 855 15607 983
rect 15676 855 15706 927
rect 15785 855 15815 927
rect 15881 855 15911 939
rect 16030 855 16060 939
rect 16121 855 16151 939
rect 16309 855 16339 985
rect 16497 855 16527 939
rect 16594 855 16624 985
<< pmos >>
rect 1814 4580 2014 4980
rect 2194 4580 2394 4980
rect 2574 4580 3574 4980
rect 3754 4580 3954 4980
rect 434 3900 634 4300
rect 814 3900 1014 4300
rect 1072 3900 1272 4300
rect 1454 3900 1654 4300
rect 1712 3900 1912 4300
rect 1970 3900 2170 4300
rect 2228 3900 2428 4300
rect 2614 3900 2814 4300
rect 2872 3900 3072 4300
rect 3130 3900 3330 4300
rect 3388 3900 3588 4300
rect 3774 3900 3974 4300
rect 414 2660 614 3060
rect 794 2660 994 3060
rect 1052 2660 1252 3060
rect 1310 2660 1510 3060
rect 1568 2660 1768 3060
rect 1826 2660 2026 3060
rect 2084 2660 2284 3060
rect 2342 2660 2542 3060
rect 2600 2660 2800 3060
rect 2974 2660 3174 3060
rect 5822 2282 6022 5282
rect 6080 2282 6280 5282
rect 6338 2282 6538 5282
rect 6596 2282 6796 5282
rect 6982 5082 7182 5282
rect 7240 5082 7440 5282
rect 7498 5082 7698 5282
rect 7756 5082 7956 5282
rect 8014 5082 8214 5282
rect 8272 5082 8472 5282
rect 8530 5082 8730 5282
rect 8902 5082 9102 5282
rect 9160 5082 9360 5282
rect 9418 5082 9618 5282
rect 9676 5082 9876 5282
rect 9934 5082 10134 5282
rect 10192 5082 10392 5282
rect 10450 5082 10650 5282
rect 10822 2282 11022 5282
rect 11080 2282 11280 5282
rect 11338 2282 11538 5282
rect 11596 2282 11796 5282
rect 17210 1153 17240 1753
<< scpmoshvt >>
rect 14677 1171 14707 1299
rect 14761 1171 14791 1299
rect 15028 1221 15058 1305
rect 15120 1221 15150 1305
rect 15219 1221 15249 1305
rect 15359 1221 15389 1305
rect 15456 1221 15486 1305
rect 15653 1137 15683 1305
rect 15752 1221 15782 1305
rect 15838 1221 15868 1305
rect 15922 1221 15952 1305
rect 16030 1221 16060 1305
rect 16114 1221 16144 1305
rect 16278 1105 16308 1305
rect 16497 1177 16527 1305
rect 16594 1105 16624 1305
<< ndiff >>
rect 8628 4598 8690 4610
rect 8628 4322 8640 4598
rect 8674 4322 8690 4598
rect 8628 4310 8690 4322
rect 8720 4598 8786 4610
rect 8720 4322 8736 4598
rect 8770 4322 8786 4598
rect 8720 4310 8786 4322
rect 8816 4598 8882 4610
rect 8816 4322 8832 4598
rect 8866 4322 8882 4598
rect 8816 4310 8882 4322
rect 8912 4598 8978 4610
rect 8912 4322 8928 4598
rect 8962 4322 8978 4598
rect 8912 4310 8978 4322
rect 9008 4598 9070 4610
rect 9008 4322 9024 4598
rect 9058 4322 9070 4598
rect 9008 4310 9070 4322
rect 7608 3878 7666 3890
rect 7608 3702 7620 3878
rect 7654 3702 7666 3878
rect 7608 3690 7666 3702
rect 7866 3878 7924 3890
rect 7866 3702 7878 3878
rect 7912 3702 7924 3878
rect 7866 3690 7924 3702
rect 8124 3878 8182 3890
rect 8124 3702 8136 3878
rect 8170 3702 8182 3878
rect 8124 3690 8182 3702
rect 8382 3878 8440 3890
rect 8382 3702 8394 3878
rect 8428 3702 8440 3878
rect 8382 3690 8440 3702
rect 8640 3878 8698 3890
rect 8640 3702 8652 3878
rect 8686 3702 8698 3878
rect 8640 3690 8698 3702
rect 8768 3818 8826 3830
rect 8768 2842 8780 3818
rect 8814 2842 8826 3818
rect 8768 2830 8826 2842
rect 9026 3818 9084 3830
rect 9026 2842 9038 3818
rect 9072 2842 9084 3818
rect 9026 2830 9084 2842
rect 9284 3818 9342 3830
rect 9284 2842 9296 3818
rect 9330 2842 9342 3818
rect 9284 2830 9342 2842
rect 9542 3818 9600 3830
rect 9542 2842 9554 3818
rect 9588 2842 9600 3818
rect 9542 2830 9600 2842
rect 9800 3818 9858 3830
rect 9800 2842 9812 3818
rect 9846 2842 9858 3818
rect 9800 2830 9858 2842
rect 10058 3818 10116 3830
rect 10058 2842 10070 3818
rect 10104 2842 10116 3818
rect 10058 2830 10116 2842
rect 10316 3818 10374 3830
rect 10316 2842 10328 3818
rect 10362 2842 10374 3818
rect 10316 2830 10374 2842
rect 160 1860 218 1872
rect 160 1684 172 1860
rect 206 1684 218 1860
rect 160 1672 218 1684
rect 418 1860 476 1872
rect 418 1684 430 1860
rect 464 1684 476 1860
rect 418 1672 476 1684
rect 540 1860 598 1872
rect 540 1684 552 1860
rect 586 1684 598 1860
rect 540 1672 598 1684
rect 798 1860 856 1872
rect 798 1684 810 1860
rect 844 1684 856 1860
rect 798 1672 856 1684
rect 920 1860 978 1872
rect 920 1684 932 1860
rect 966 1684 978 1860
rect 920 1672 978 1684
rect 1178 1860 1236 1872
rect 1178 1684 1190 1860
rect 1224 1684 1236 1860
rect 1178 1672 1236 1684
rect 1300 1860 1358 1872
rect 1300 1684 1312 1860
rect 1346 1684 1358 1860
rect 1300 1672 1358 1684
rect 1558 1860 1616 1872
rect 1558 1684 1570 1860
rect 1604 1684 1616 1860
rect 1558 1672 1616 1684
rect 1680 1860 1738 1872
rect 1680 1684 1692 1860
rect 1726 1684 1738 1860
rect 1680 1672 1738 1684
rect 1938 1860 1996 1872
rect 1938 1684 1950 1860
rect 1984 1684 1996 1860
rect 1938 1672 1996 1684
rect 2060 1860 2118 1872
rect 2060 1684 2072 1860
rect 2106 1684 2118 1860
rect 2060 1672 2118 1684
rect 2318 1860 2376 1872
rect 2318 1684 2330 1860
rect 2364 1684 2376 1860
rect 2318 1672 2376 1684
rect 2440 1860 2498 1872
rect 2440 1684 2452 1860
rect 2486 1684 2498 1860
rect 2440 1672 2498 1684
rect 2698 1860 2756 1872
rect 2698 1684 2710 1860
rect 2744 1684 2756 1860
rect 2698 1672 2756 1684
rect 2820 1860 2878 1872
rect 2820 1684 2832 1860
rect 2866 1684 2878 1860
rect 2820 1672 2878 1684
rect 3078 1860 3136 1872
rect 3078 1684 3090 1860
rect 3124 1684 3136 1860
rect 3078 1672 3136 1684
rect 160 1442 218 1454
rect 160 1266 172 1442
rect 206 1266 218 1442
rect 160 1254 218 1266
rect 418 1442 476 1454
rect 418 1266 430 1442
rect 464 1266 476 1442
rect 418 1254 476 1266
rect 540 1442 598 1454
rect 540 1266 552 1442
rect 586 1266 598 1442
rect 540 1254 598 1266
rect 798 1442 856 1454
rect 798 1266 810 1442
rect 844 1266 856 1442
rect 798 1254 856 1266
rect 920 1442 978 1454
rect 920 1266 932 1442
rect 966 1266 978 1442
rect 920 1254 978 1266
rect 1178 1442 1236 1454
rect 1178 1266 1190 1442
rect 1224 1266 1236 1442
rect 1178 1254 1236 1266
rect 1300 1442 1358 1454
rect 1300 1266 1312 1442
rect 1346 1266 1358 1442
rect 1300 1254 1358 1266
rect 1558 1442 1616 1454
rect 1558 1266 1570 1442
rect 1604 1266 1616 1442
rect 1558 1254 1616 1266
rect 1680 1442 1738 1454
rect 1680 1266 1692 1442
rect 1726 1266 1738 1442
rect 1680 1254 1738 1266
rect 1938 1442 1996 1454
rect 1938 1266 1950 1442
rect 1984 1266 1996 1442
rect 1938 1254 1996 1266
rect 2060 1442 2118 1454
rect 2060 1266 2072 1442
rect 2106 1266 2118 1442
rect 2060 1254 2118 1266
rect 2318 1442 2376 1454
rect 2318 1266 2330 1442
rect 2364 1266 2376 1442
rect 2318 1254 2376 1266
rect 2440 1442 2498 1454
rect 2440 1266 2452 1442
rect 2486 1266 2498 1442
rect 2440 1254 2498 1266
rect 2698 1442 2756 1454
rect 2698 1266 2710 1442
rect 2744 1266 2756 1442
rect 2698 1254 2756 1266
rect 2820 1442 2878 1454
rect 2820 1266 2832 1442
rect 2866 1266 2878 1442
rect 2820 1254 2878 1266
rect 3078 1442 3136 1454
rect 3078 1266 3090 1442
rect 3124 1266 3136 1442
rect 3078 1254 3136 1266
rect 160 1024 218 1036
rect 160 848 172 1024
rect 206 848 218 1024
rect 160 836 218 848
rect 418 1024 476 1036
rect 418 848 430 1024
rect 464 848 476 1024
rect 418 836 476 848
rect 540 1024 598 1036
rect 540 848 552 1024
rect 586 848 598 1024
rect 540 836 598 848
rect 798 1024 856 1036
rect 798 848 810 1024
rect 844 848 856 1024
rect 798 836 856 848
rect 920 1024 978 1036
rect 920 848 932 1024
rect 966 848 978 1024
rect 920 836 978 848
rect 1178 1024 1236 1036
rect 1178 848 1190 1024
rect 1224 848 1236 1024
rect 1178 836 1236 848
rect 1300 1024 1358 1036
rect 1300 848 1312 1024
rect 1346 848 1358 1024
rect 1300 836 1358 848
rect 1558 1024 1616 1036
rect 1558 848 1570 1024
rect 1604 848 1616 1024
rect 1558 836 1616 848
rect 1680 1024 1738 1036
rect 1680 848 1692 1024
rect 1726 848 1738 1024
rect 1680 836 1738 848
rect 1938 1024 1996 1036
rect 1938 848 1950 1024
rect 1984 848 1996 1024
rect 1938 836 1996 848
rect 2060 1024 2118 1036
rect 2060 848 2072 1024
rect 2106 848 2118 1024
rect 2060 836 2118 848
rect 2318 1024 2376 1036
rect 2318 848 2330 1024
rect 2364 848 2376 1024
rect 2318 836 2376 848
rect 2440 1024 2498 1036
rect 2440 848 2452 1024
rect 2486 848 2498 1024
rect 2440 836 2498 848
rect 2698 1024 2756 1036
rect 2698 848 2710 1024
rect 2744 848 2756 1024
rect 2698 836 2756 848
rect 2820 1024 2878 1036
rect 2820 848 2832 1024
rect 2866 848 2878 1024
rect 2820 836 2878 848
rect 3078 1024 3136 1036
rect 3078 848 3090 1024
rect 3124 848 3136 1024
rect 3078 836 3136 848
rect 160 606 218 618
rect 160 430 172 606
rect 206 430 218 606
rect 160 418 218 430
rect 418 606 476 618
rect 418 430 430 606
rect 464 430 476 606
rect 418 418 476 430
rect 540 606 598 618
rect 540 430 552 606
rect 586 430 598 606
rect 540 418 598 430
rect 798 606 856 618
rect 798 430 810 606
rect 844 430 856 606
rect 798 418 856 430
rect 920 606 978 618
rect 920 430 932 606
rect 966 430 978 606
rect 920 418 978 430
rect 1178 606 1236 618
rect 1178 430 1190 606
rect 1224 430 1236 606
rect 1178 418 1236 430
rect 1300 606 1358 618
rect 1300 430 1312 606
rect 1346 430 1358 606
rect 1300 418 1358 430
rect 1558 606 1616 618
rect 1558 430 1570 606
rect 1604 430 1616 606
rect 1558 418 1616 430
rect 1680 606 1738 618
rect 1680 430 1692 606
rect 1726 430 1738 606
rect 1680 418 1738 430
rect 1938 606 1996 618
rect 1938 430 1950 606
rect 1984 430 1996 606
rect 1938 418 1996 430
rect 2060 606 2118 618
rect 2060 430 2072 606
rect 2106 430 2118 606
rect 2060 418 2118 430
rect 2318 606 2376 618
rect 2318 430 2330 606
rect 2364 430 2376 606
rect 2318 418 2376 430
rect 2440 606 2498 618
rect 2440 430 2452 606
rect 2486 430 2498 606
rect 2440 418 2498 430
rect 2698 606 2756 618
rect 2698 430 2710 606
rect 2744 430 2756 606
rect 2698 418 2756 430
rect 2820 606 2878 618
rect 2820 430 2832 606
rect 2866 430 2878 606
rect 2820 418 2878 430
rect 3078 606 3136 618
rect 3078 430 3090 606
rect 3124 430 3136 606
rect 3078 418 3136 430
rect 14625 927 14677 939
rect 14625 893 14633 927
rect 14667 893 14677 927
rect 14625 855 14677 893
rect 14707 901 14761 939
rect 14707 867 14717 901
rect 14751 867 14761 901
rect 14707 855 14761 867
rect 14791 927 14843 939
rect 14791 893 14801 927
rect 14835 893 14843 927
rect 14791 855 14843 893
rect 14911 897 15016 939
rect 14911 863 14923 897
rect 14957 863 15016 897
rect 14911 855 15016 863
rect 15046 927 15096 939
rect 15527 939 15577 983
rect 15255 927 15373 939
rect 15046 903 15111 927
rect 15046 869 15056 903
rect 15090 869 15111 903
rect 15046 855 15111 869
rect 15141 903 15207 927
rect 15141 869 15163 903
rect 15197 869 15207 903
rect 15141 855 15207 869
rect 15237 855 15373 927
rect 15403 855 15445 939
rect 15475 901 15577 939
rect 15475 867 15509 901
rect 15543 867 15577 901
rect 15475 855 15577 867
rect 15607 927 15661 983
rect 16257 940 16309 985
rect 15831 927 15881 939
rect 15607 897 15676 927
rect 15607 863 15621 897
rect 15655 863 15676 897
rect 15607 855 15676 863
rect 15706 901 15785 927
rect 15706 867 15731 901
rect 15765 867 15785 901
rect 15706 855 15785 867
rect 15815 855 15881 927
rect 15911 897 16030 939
rect 15911 863 15943 897
rect 15977 863 16030 897
rect 15911 855 16030 863
rect 16060 855 16121 939
rect 16151 917 16203 939
rect 16151 883 16161 917
rect 16195 883 16203 917
rect 16151 855 16203 883
rect 16257 906 16265 940
rect 16299 906 16309 940
rect 16257 855 16309 906
rect 16339 973 16391 985
rect 16339 939 16349 973
rect 16383 939 16391 973
rect 16542 939 16594 985
rect 16339 905 16391 939
rect 16339 871 16349 905
rect 16383 871 16391 905
rect 16339 855 16391 871
rect 16445 927 16497 939
rect 16445 893 16453 927
rect 16487 893 16497 927
rect 16445 855 16497 893
rect 16527 921 16594 939
rect 16527 887 16550 921
rect 16584 887 16594 921
rect 16527 855 16594 887
rect 16624 951 16676 985
rect 16624 917 16634 951
rect 16668 917 16676 951
rect 16624 855 16676 917
rect 17152 662 17210 674
rect 17152 486 17164 662
rect 17198 486 17210 662
rect 17152 474 17210 486
rect 17240 662 17298 674
rect 17240 486 17252 662
rect 17286 486 17298 662
rect 17240 474 17298 486
<< pdiff >>
rect 1756 4968 1814 4980
rect 1756 4592 1768 4968
rect 1802 4592 1814 4968
rect 1756 4580 1814 4592
rect 2014 4968 2072 4980
rect 2014 4592 2026 4968
rect 2060 4592 2072 4968
rect 2014 4580 2072 4592
rect 2136 4968 2194 4980
rect 2136 4592 2148 4968
rect 2182 4592 2194 4968
rect 2136 4580 2194 4592
rect 2394 4968 2452 4980
rect 2394 4592 2406 4968
rect 2440 4592 2452 4968
rect 2394 4580 2452 4592
rect 2516 4968 2574 4980
rect 2516 4592 2528 4968
rect 2562 4592 2574 4968
rect 2516 4580 2574 4592
rect 3574 4968 3632 4980
rect 3574 4592 3586 4968
rect 3620 4592 3632 4968
rect 3574 4580 3632 4592
rect 3696 4968 3754 4980
rect 3696 4592 3708 4968
rect 3742 4592 3754 4968
rect 3696 4580 3754 4592
rect 3954 4968 4012 4980
rect 3954 4592 3966 4968
rect 4000 4592 4012 4968
rect 3954 4580 4012 4592
rect 376 4288 434 4300
rect 376 3912 388 4288
rect 422 3912 434 4288
rect 376 3900 434 3912
rect 634 4288 692 4300
rect 634 3912 646 4288
rect 680 3912 692 4288
rect 634 3900 692 3912
rect 756 4288 814 4300
rect 756 3912 768 4288
rect 802 3912 814 4288
rect 756 3900 814 3912
rect 1014 4288 1072 4300
rect 1014 3912 1026 4288
rect 1060 3912 1072 4288
rect 1014 3900 1072 3912
rect 1272 4288 1330 4300
rect 1272 3912 1284 4288
rect 1318 3912 1330 4288
rect 1272 3900 1330 3912
rect 1396 4288 1454 4300
rect 1396 3912 1408 4288
rect 1442 3912 1454 4288
rect 1396 3900 1454 3912
rect 1654 4288 1712 4300
rect 1654 3912 1666 4288
rect 1700 3912 1712 4288
rect 1654 3900 1712 3912
rect 1912 4288 1970 4300
rect 1912 3912 1924 4288
rect 1958 3912 1970 4288
rect 1912 3900 1970 3912
rect 2170 4288 2228 4300
rect 2170 3912 2182 4288
rect 2216 3912 2228 4288
rect 2170 3900 2228 3912
rect 2428 4288 2486 4300
rect 2428 3912 2440 4288
rect 2474 3912 2486 4288
rect 2428 3900 2486 3912
rect 2556 4288 2614 4300
rect 2556 3912 2568 4288
rect 2602 3912 2614 4288
rect 2556 3900 2614 3912
rect 2814 4288 2872 4300
rect 2814 3912 2826 4288
rect 2860 3912 2872 4288
rect 2814 3900 2872 3912
rect 3072 4288 3130 4300
rect 3072 3912 3084 4288
rect 3118 3912 3130 4288
rect 3072 3900 3130 3912
rect 3330 4288 3388 4300
rect 3330 3912 3342 4288
rect 3376 3912 3388 4288
rect 3330 3900 3388 3912
rect 3588 4288 3646 4300
rect 3588 3912 3600 4288
rect 3634 3912 3646 4288
rect 3588 3900 3646 3912
rect 3716 4288 3774 4300
rect 3716 3912 3728 4288
rect 3762 3912 3774 4288
rect 3716 3900 3774 3912
rect 3974 4288 4032 4300
rect 3974 3912 3986 4288
rect 4020 3912 4032 4288
rect 3974 3900 4032 3912
rect 356 3048 414 3060
rect 356 2672 368 3048
rect 402 2672 414 3048
rect 356 2660 414 2672
rect 614 3048 672 3060
rect 614 2672 626 3048
rect 660 2672 672 3048
rect 614 2660 672 2672
rect 736 3048 794 3060
rect 736 2672 748 3048
rect 782 2672 794 3048
rect 736 2660 794 2672
rect 994 3048 1052 3060
rect 994 2672 1006 3048
rect 1040 2672 1052 3048
rect 994 2660 1052 2672
rect 1252 3048 1310 3060
rect 1252 2672 1264 3048
rect 1298 2672 1310 3048
rect 1252 2660 1310 2672
rect 1510 3048 1568 3060
rect 1510 2672 1522 3048
rect 1556 2672 1568 3048
rect 1510 2660 1568 2672
rect 1768 3048 1826 3060
rect 1768 2672 1780 3048
rect 1814 2672 1826 3048
rect 1768 2660 1826 2672
rect 2026 3048 2084 3060
rect 2026 2672 2038 3048
rect 2072 2672 2084 3048
rect 2026 2660 2084 2672
rect 2284 3048 2342 3060
rect 2284 2672 2296 3048
rect 2330 2672 2342 3048
rect 2284 2660 2342 2672
rect 2542 3048 2600 3060
rect 2542 2672 2554 3048
rect 2588 2672 2600 3048
rect 2542 2660 2600 2672
rect 2800 3048 2858 3060
rect 2800 2672 2812 3048
rect 2846 2672 2858 3048
rect 2800 2660 2858 2672
rect 2916 3048 2974 3060
rect 2916 2672 2928 3048
rect 2962 2672 2974 3048
rect 2916 2660 2974 2672
rect 3174 3048 3232 3060
rect 3174 2672 3186 3048
rect 3220 2672 3232 3048
rect 3174 2660 3232 2672
rect 5764 5270 5822 5282
rect 5764 2294 5776 5270
rect 5810 2294 5822 5270
rect 5764 2282 5822 2294
rect 6022 5270 6080 5282
rect 6022 2294 6034 5270
rect 6068 2294 6080 5270
rect 6022 2282 6080 2294
rect 6280 5270 6338 5282
rect 6280 2294 6292 5270
rect 6326 2294 6338 5270
rect 6280 2282 6338 2294
rect 6538 5270 6596 5282
rect 6538 2294 6550 5270
rect 6584 2294 6596 5270
rect 6538 2282 6596 2294
rect 6796 5270 6854 5282
rect 6796 2294 6808 5270
rect 6842 2294 6854 5270
rect 6924 5270 6982 5282
rect 6924 5094 6936 5270
rect 6970 5094 6982 5270
rect 6924 5082 6982 5094
rect 7182 5270 7240 5282
rect 7182 5094 7194 5270
rect 7228 5094 7240 5270
rect 7182 5082 7240 5094
rect 7440 5270 7498 5282
rect 7440 5094 7452 5270
rect 7486 5094 7498 5270
rect 7440 5082 7498 5094
rect 7698 5270 7756 5282
rect 7698 5094 7710 5270
rect 7744 5094 7756 5270
rect 7698 5082 7756 5094
rect 7956 5270 8014 5282
rect 7956 5094 7968 5270
rect 8002 5094 8014 5270
rect 7956 5082 8014 5094
rect 8214 5270 8272 5282
rect 8214 5094 8226 5270
rect 8260 5094 8272 5270
rect 8214 5082 8272 5094
rect 8472 5270 8530 5282
rect 8472 5094 8484 5270
rect 8518 5094 8530 5270
rect 8472 5082 8530 5094
rect 8730 5270 8788 5282
rect 8730 5094 8742 5270
rect 8776 5094 8788 5270
rect 8730 5082 8788 5094
rect 8844 5270 8902 5282
rect 8844 5094 8856 5270
rect 8890 5094 8902 5270
rect 8844 5082 8902 5094
rect 9102 5270 9160 5282
rect 9102 5094 9114 5270
rect 9148 5094 9160 5270
rect 9102 5082 9160 5094
rect 9360 5270 9418 5282
rect 9360 5094 9372 5270
rect 9406 5094 9418 5270
rect 9360 5082 9418 5094
rect 9618 5270 9676 5282
rect 9618 5094 9630 5270
rect 9664 5094 9676 5270
rect 9618 5082 9676 5094
rect 9876 5270 9934 5282
rect 9876 5094 9888 5270
rect 9922 5094 9934 5270
rect 9876 5082 9934 5094
rect 10134 5270 10192 5282
rect 10134 5094 10146 5270
rect 10180 5094 10192 5270
rect 10134 5082 10192 5094
rect 10392 5270 10450 5282
rect 10392 5094 10404 5270
rect 10438 5094 10450 5270
rect 10392 5082 10450 5094
rect 10650 5270 10708 5282
rect 10650 5094 10662 5270
rect 10696 5094 10708 5270
rect 10650 5082 10708 5094
rect 10764 5270 10822 5282
rect 6796 2282 6854 2294
rect 10764 2294 10776 5270
rect 10810 2294 10822 5270
rect 10764 2282 10822 2294
rect 11022 5270 11080 5282
rect 11022 2294 11034 5270
rect 11068 2294 11080 5270
rect 11022 2282 11080 2294
rect 11280 5270 11338 5282
rect 11280 2294 11292 5270
rect 11326 2294 11338 5270
rect 11280 2282 11338 2294
rect 11538 5270 11596 5282
rect 11538 2294 11550 5270
rect 11584 2294 11596 5270
rect 11538 2282 11596 2294
rect 11796 5270 11854 5282
rect 11796 2294 11808 5270
rect 11842 2294 11854 5270
rect 11796 2282 11854 2294
rect 14625 1285 14677 1299
rect 14625 1251 14633 1285
rect 14667 1251 14677 1285
rect 14625 1217 14677 1251
rect 14625 1183 14633 1217
rect 14667 1183 14677 1217
rect 14625 1171 14677 1183
rect 14707 1269 14761 1299
rect 14707 1235 14717 1269
rect 14751 1235 14761 1269
rect 14707 1171 14761 1235
rect 14791 1285 14843 1299
rect 14791 1251 14801 1285
rect 14835 1251 14843 1285
rect 14791 1217 14843 1251
rect 14976 1293 15028 1305
rect 14976 1259 14984 1293
rect 15018 1259 15028 1293
rect 14976 1221 15028 1259
rect 15058 1285 15120 1305
rect 15058 1251 15068 1285
rect 15102 1251 15120 1285
rect 15058 1221 15120 1251
rect 15150 1291 15219 1305
rect 15150 1257 15161 1291
rect 15195 1257 15219 1291
rect 15150 1221 15219 1257
rect 15249 1267 15359 1305
rect 15249 1233 15315 1267
rect 15349 1233 15359 1267
rect 15249 1221 15359 1233
rect 15389 1283 15456 1305
rect 15389 1249 15412 1283
rect 15446 1249 15456 1283
rect 15389 1221 15456 1249
rect 15486 1267 15538 1305
rect 15486 1233 15496 1267
rect 15530 1233 15538 1267
rect 15486 1221 15538 1233
rect 15601 1293 15653 1305
rect 15601 1259 15609 1293
rect 15643 1259 15653 1293
rect 14791 1183 14801 1217
rect 14835 1183 14843 1217
rect 14791 1171 14843 1183
rect 15601 1137 15653 1259
rect 15683 1285 15752 1305
rect 15683 1251 15697 1285
rect 15731 1251 15752 1285
rect 15683 1221 15752 1251
rect 15782 1292 15838 1305
rect 15782 1258 15794 1292
rect 15828 1258 15838 1292
rect 15782 1221 15838 1258
rect 15868 1221 15922 1305
rect 15952 1293 16030 1305
rect 15952 1259 15986 1293
rect 16020 1259 16030 1293
rect 15952 1221 16030 1259
rect 16060 1267 16114 1305
rect 16060 1233 16070 1267
rect 16104 1233 16114 1267
rect 16060 1221 16114 1233
rect 16144 1293 16278 1305
rect 16144 1259 16156 1293
rect 16190 1259 16234 1293
rect 16268 1259 16278 1293
rect 16144 1221 16278 1259
rect 15683 1137 15737 1221
rect 16228 1105 16278 1221
rect 16308 1285 16364 1305
rect 16308 1251 16318 1285
rect 16352 1251 16364 1285
rect 16308 1217 16364 1251
rect 16308 1183 16318 1217
rect 16352 1183 16364 1217
rect 16308 1149 16364 1183
rect 16445 1293 16497 1305
rect 16445 1259 16453 1293
rect 16487 1259 16497 1293
rect 16445 1225 16497 1259
rect 16445 1191 16453 1225
rect 16487 1191 16497 1225
rect 16445 1177 16497 1191
rect 16527 1293 16594 1305
rect 16527 1259 16550 1293
rect 16584 1259 16594 1293
rect 16527 1225 16594 1259
rect 16527 1191 16550 1225
rect 16584 1191 16594 1225
rect 16527 1177 16594 1191
rect 16308 1115 16318 1149
rect 16352 1115 16364 1149
rect 16308 1105 16364 1115
rect 16542 1157 16594 1177
rect 16542 1123 16550 1157
rect 16584 1123 16594 1157
rect 16542 1105 16594 1123
rect 16624 1257 16676 1305
rect 16624 1223 16634 1257
rect 16668 1223 16676 1257
rect 16624 1189 16676 1223
rect 16624 1155 16634 1189
rect 16668 1155 16676 1189
rect 16624 1105 16676 1155
rect 17152 1741 17210 1753
rect 17152 1165 17164 1741
rect 17198 1165 17210 1741
rect 17152 1153 17210 1165
rect 17240 1741 17298 1753
rect 17240 1165 17252 1741
rect 17286 1165 17298 1741
rect 17240 1153 17298 1165
<< ndiffc >>
rect 8640 4322 8674 4598
rect 8736 4322 8770 4598
rect 8832 4322 8866 4598
rect 8928 4322 8962 4598
rect 9024 4322 9058 4598
rect 7620 3702 7654 3878
rect 7878 3702 7912 3878
rect 8136 3702 8170 3878
rect 8394 3702 8428 3878
rect 8652 3702 8686 3878
rect 8780 2842 8814 3818
rect 9038 2842 9072 3818
rect 9296 2842 9330 3818
rect 9554 2842 9588 3818
rect 9812 2842 9846 3818
rect 10070 2842 10104 3818
rect 10328 2842 10362 3818
rect 172 1684 206 1860
rect 430 1684 464 1860
rect 552 1684 586 1860
rect 810 1684 844 1860
rect 932 1684 966 1860
rect 1190 1684 1224 1860
rect 1312 1684 1346 1860
rect 1570 1684 1604 1860
rect 1692 1684 1726 1860
rect 1950 1684 1984 1860
rect 2072 1684 2106 1860
rect 2330 1684 2364 1860
rect 2452 1684 2486 1860
rect 2710 1684 2744 1860
rect 2832 1684 2866 1860
rect 3090 1684 3124 1860
rect 172 1266 206 1442
rect 430 1266 464 1442
rect 552 1266 586 1442
rect 810 1266 844 1442
rect 932 1266 966 1442
rect 1190 1266 1224 1442
rect 1312 1266 1346 1442
rect 1570 1266 1604 1442
rect 1692 1266 1726 1442
rect 1950 1266 1984 1442
rect 2072 1266 2106 1442
rect 2330 1266 2364 1442
rect 2452 1266 2486 1442
rect 2710 1266 2744 1442
rect 2832 1266 2866 1442
rect 3090 1266 3124 1442
rect 172 848 206 1024
rect 430 848 464 1024
rect 552 848 586 1024
rect 810 848 844 1024
rect 932 848 966 1024
rect 1190 848 1224 1024
rect 1312 848 1346 1024
rect 1570 848 1604 1024
rect 1692 848 1726 1024
rect 1950 848 1984 1024
rect 2072 848 2106 1024
rect 2330 848 2364 1024
rect 2452 848 2486 1024
rect 2710 848 2744 1024
rect 2832 848 2866 1024
rect 3090 848 3124 1024
rect 172 430 206 606
rect 430 430 464 606
rect 552 430 586 606
rect 810 430 844 606
rect 932 430 966 606
rect 1190 430 1224 606
rect 1312 430 1346 606
rect 1570 430 1604 606
rect 1692 430 1726 606
rect 1950 430 1984 606
rect 2072 430 2106 606
rect 2330 430 2364 606
rect 2452 430 2486 606
rect 2710 430 2744 606
rect 2832 430 2866 606
rect 3090 430 3124 606
rect 14633 893 14667 927
rect 14717 867 14751 901
rect 14801 893 14835 927
rect 14923 863 14957 897
rect 15056 869 15090 903
rect 15163 869 15197 903
rect 15509 867 15543 901
rect 15621 863 15655 897
rect 15731 867 15765 901
rect 15943 863 15977 897
rect 16161 883 16195 917
rect 16265 906 16299 940
rect 16349 939 16383 973
rect 16349 871 16383 905
rect 16453 893 16487 927
rect 16550 887 16584 921
rect 16634 917 16668 951
rect 17164 486 17198 662
rect 17252 486 17286 662
<< pdiffc >>
rect 1768 4592 1802 4968
rect 2026 4592 2060 4968
rect 2148 4592 2182 4968
rect 2406 4592 2440 4968
rect 2528 4592 2562 4968
rect 3586 4592 3620 4968
rect 3708 4592 3742 4968
rect 3966 4592 4000 4968
rect 388 3912 422 4288
rect 646 3912 680 4288
rect 768 3912 802 4288
rect 1026 3912 1060 4288
rect 1284 3912 1318 4288
rect 1408 3912 1442 4288
rect 1666 3912 1700 4288
rect 1924 3912 1958 4288
rect 2182 3912 2216 4288
rect 2440 3912 2474 4288
rect 2568 3912 2602 4288
rect 2826 3912 2860 4288
rect 3084 3912 3118 4288
rect 3342 3912 3376 4288
rect 3600 3912 3634 4288
rect 3728 3912 3762 4288
rect 3986 3912 4020 4288
rect 368 2672 402 3048
rect 626 2672 660 3048
rect 748 2672 782 3048
rect 1006 2672 1040 3048
rect 1264 2672 1298 3048
rect 1522 2672 1556 3048
rect 1780 2672 1814 3048
rect 2038 2672 2072 3048
rect 2296 2672 2330 3048
rect 2554 2672 2588 3048
rect 2812 2672 2846 3048
rect 2928 2672 2962 3048
rect 3186 2672 3220 3048
rect 5776 2294 5810 5270
rect 6034 2294 6068 5270
rect 6292 2294 6326 5270
rect 6550 2294 6584 5270
rect 6808 2294 6842 5270
rect 6936 5094 6970 5270
rect 7194 5094 7228 5270
rect 7452 5094 7486 5270
rect 7710 5094 7744 5270
rect 7968 5094 8002 5270
rect 8226 5094 8260 5270
rect 8484 5094 8518 5270
rect 8742 5094 8776 5270
rect 8856 5094 8890 5270
rect 9114 5094 9148 5270
rect 9372 5094 9406 5270
rect 9630 5094 9664 5270
rect 9888 5094 9922 5270
rect 10146 5094 10180 5270
rect 10404 5094 10438 5270
rect 10662 5094 10696 5270
rect 10776 2294 10810 5270
rect 11034 2294 11068 5270
rect 11292 2294 11326 5270
rect 11550 2294 11584 5270
rect 11808 2294 11842 5270
rect 14633 1251 14667 1285
rect 14633 1183 14667 1217
rect 14717 1235 14751 1269
rect 14801 1251 14835 1285
rect 14984 1259 15018 1293
rect 15068 1251 15102 1285
rect 15161 1257 15195 1291
rect 15315 1233 15349 1267
rect 15412 1249 15446 1283
rect 15496 1233 15530 1267
rect 15609 1259 15643 1293
rect 14801 1183 14835 1217
rect 15697 1251 15731 1285
rect 15794 1258 15828 1292
rect 15986 1259 16020 1293
rect 16070 1233 16104 1267
rect 16156 1259 16190 1293
rect 16234 1259 16268 1293
rect 16318 1251 16352 1285
rect 16318 1183 16352 1217
rect 16453 1259 16487 1293
rect 16453 1191 16487 1225
rect 16550 1259 16584 1293
rect 16550 1191 16584 1225
rect 16318 1115 16352 1149
rect 16550 1123 16584 1157
rect 16634 1223 16668 1257
rect 16634 1155 16668 1189
rect 17164 1165 17198 1741
rect 17252 1165 17286 1741
<< psubdiff >>
rect 14396 5870 14492 5904
rect 17420 5870 17516 5904
rect 14396 5808 14430 5870
rect 7344 4732 7440 4766
rect 10368 4732 10464 4766
rect 7344 4670 7378 4732
rect 10430 4670 10464 4732
rect 7344 2652 7378 2714
rect 10430 2652 10464 2714
rect 7344 2618 7440 2652
rect 10368 2618 10464 2652
rect 17482 5808 17516 5870
rect 14396 2190 14430 2252
rect 17482 2190 17516 2252
rect 14396 2156 14492 2190
rect 17420 2156 17516 2190
rect 36 2010 132 2044
rect 3260 2010 3356 2044
rect 36 1948 70 2010
rect 3322 1948 3356 2010
rect 36 230 70 292
rect 17050 814 17146 848
rect 17304 814 17400 848
rect 17050 752 17084 814
rect 17366 752 17400 814
rect 17050 334 17084 396
rect 17366 334 17400 396
rect 17050 300 17146 334
rect 17304 300 17400 334
rect 3322 230 3356 292
rect 36 196 132 230
rect 3260 196 3356 230
<< nsubdiff >>
rect 11848 5499 11948 5502
rect 5671 5465 5731 5499
rect 11885 5465 11948 5499
rect 5671 5439 5705 5465
rect 7071 5462 7105 5465
rect 10571 5462 10605 5465
rect 11848 5462 11948 5465
rect 243 5223 303 5257
rect 4137 5223 4197 5257
rect 243 5197 277 5223
rect 4163 5197 4197 5223
rect 243 3697 277 3723
rect 4163 3697 4197 3723
rect 243 3663 303 3697
rect 4137 3663 4197 3697
rect 203 3303 263 3337
rect 3297 3303 3357 3337
rect 203 3277 237 3303
rect 3323 3277 3357 3303
rect 203 2377 237 2403
rect 3323 2377 3357 2403
rect 203 2343 263 2377
rect 3297 2343 3357 2377
rect 11911 5439 11945 5462
rect 5705 4845 5708 4879
rect 6948 4879 7208 4882
rect 10671 4879 10705 4882
rect 6928 4845 7148 4879
rect 10528 4845 10705 4879
rect 6928 4842 7208 4845
rect 6928 4765 6965 4842
rect 10671 4802 10705 4845
rect 6931 4762 6965 4765
rect 5671 2119 5705 2145
rect 6931 2119 6965 2145
rect 5671 2085 5731 2119
rect 6905 2085 6965 2119
rect 11908 4845 11911 4879
rect 10671 2119 10705 2145
rect 11911 2119 11945 2145
rect 10671 2085 10731 2119
rect 11885 2085 11945 2119
rect 17050 1902 17146 1936
rect 17304 1902 17400 1936
rect 17050 1840 17084 1902
rect 14420 1290 14520 1310
rect 14420 1250 14450 1290
rect 14490 1250 14520 1290
rect 14420 1220 14520 1250
rect 17366 1840 17400 1902
rect 17050 1004 17084 1066
rect 17366 1004 17400 1066
rect 17050 970 17146 1004
rect 17304 970 17400 1004
<< psubdiffcont >>
rect 14492 5870 17420 5904
rect 7440 4732 10368 4766
rect 7344 2714 7378 4670
rect 10430 2714 10464 4670
rect 7440 2618 10368 2652
rect 14396 2252 14430 5808
rect 17482 2252 17516 5808
rect 14492 2156 17420 2190
rect 132 2010 3260 2044
rect 36 292 70 1948
rect 3322 292 3356 1948
rect 17146 814 17304 848
rect 17050 396 17084 752
rect 17366 396 17400 752
rect 17146 300 17304 334
rect 132 196 3260 230
<< nsubdiffcont >>
rect 5731 5465 11885 5499
rect 303 5223 4137 5257
rect 243 3723 277 5197
rect 4163 3723 4197 5197
rect 303 3663 4137 3697
rect 263 3303 3297 3337
rect 203 2403 237 3277
rect 3323 2403 3357 3277
rect 263 2343 3297 2377
rect 5671 2145 5705 5439
rect 7148 4845 10528 4879
rect 6931 2145 6965 4762
rect 5731 2085 6905 2119
rect 10671 2145 10705 4802
rect 11911 2145 11945 5439
rect 10731 2085 11885 2119
rect 17146 1902 17304 1936
rect 14450 1250 14490 1290
rect 17050 1066 17084 1840
rect 17366 1066 17400 1840
rect 17146 970 17304 1004
<< poly >>
rect 1814 5061 2014 5077
rect 1814 5027 1830 5061
rect 1998 5027 2014 5061
rect 1814 4980 2014 5027
rect 2194 5061 2394 5077
rect 2194 5027 2210 5061
rect 2378 5027 2394 5061
rect 2194 4980 2394 5027
rect 2574 5061 3574 5077
rect 2574 5027 2590 5061
rect 3558 5027 3574 5061
rect 2574 4980 3574 5027
rect 3754 5061 3954 5077
rect 3754 5027 3770 5061
rect 3938 5027 3954 5061
rect 3754 4980 3954 5027
rect 1814 4533 2014 4580
rect 1814 4499 1830 4533
rect 1998 4499 2014 4533
rect 1814 4483 2014 4499
rect 2194 4533 2394 4580
rect 2194 4499 2210 4533
rect 2378 4499 2394 4533
rect 2194 4483 2394 4499
rect 2574 4533 3574 4580
rect 2574 4499 2590 4533
rect 3558 4499 3574 4533
rect 2574 4483 3574 4499
rect 3754 4533 3954 4580
rect 3754 4499 3770 4533
rect 3938 4499 3954 4533
rect 3754 4483 3954 4499
rect 434 4381 634 4397
rect 434 4347 450 4381
rect 618 4347 634 4381
rect 434 4300 634 4347
rect 814 4381 1014 4397
rect 814 4347 830 4381
rect 998 4347 1014 4381
rect 814 4300 1014 4347
rect 1072 4381 1272 4397
rect 1072 4347 1088 4381
rect 1256 4347 1272 4381
rect 1072 4300 1272 4347
rect 1454 4381 1654 4397
rect 1454 4347 1470 4381
rect 1638 4347 1654 4381
rect 1454 4300 1654 4347
rect 1712 4381 1912 4397
rect 1712 4347 1728 4381
rect 1896 4347 1912 4381
rect 1712 4300 1912 4347
rect 1970 4381 2170 4397
rect 1970 4347 1986 4381
rect 2154 4347 2170 4381
rect 1970 4300 2170 4347
rect 2228 4381 2428 4397
rect 2228 4347 2244 4381
rect 2412 4347 2428 4381
rect 2228 4300 2428 4347
rect 2614 4381 2814 4397
rect 2614 4347 2630 4381
rect 2798 4347 2814 4381
rect 2614 4300 2814 4347
rect 2872 4381 3072 4397
rect 2872 4347 2888 4381
rect 3056 4347 3072 4381
rect 2872 4300 3072 4347
rect 3130 4381 3330 4397
rect 3130 4347 3146 4381
rect 3314 4347 3330 4381
rect 3130 4300 3330 4347
rect 3388 4381 3588 4397
rect 3388 4347 3404 4381
rect 3572 4347 3588 4381
rect 3388 4300 3588 4347
rect 3774 4381 3974 4397
rect 3774 4347 3790 4381
rect 3958 4347 3974 4381
rect 3774 4300 3974 4347
rect 434 3853 634 3900
rect 434 3819 450 3853
rect 618 3819 634 3853
rect 434 3803 634 3819
rect 814 3853 1014 3900
rect 814 3819 830 3853
rect 998 3819 1014 3853
rect 814 3803 1014 3819
rect 1072 3853 1272 3900
rect 1072 3819 1088 3853
rect 1256 3819 1272 3853
rect 1072 3803 1272 3819
rect 1454 3853 1654 3900
rect 1454 3819 1470 3853
rect 1638 3819 1654 3853
rect 1454 3803 1654 3819
rect 1712 3853 1912 3900
rect 1712 3819 1728 3853
rect 1896 3819 1912 3853
rect 1712 3803 1912 3819
rect 1970 3853 2170 3900
rect 1970 3819 1986 3853
rect 2154 3819 2170 3853
rect 1970 3803 2170 3819
rect 2228 3853 2428 3900
rect 2228 3819 2244 3853
rect 2412 3819 2428 3853
rect 2228 3803 2428 3819
rect 2614 3853 2814 3900
rect 2614 3819 2630 3853
rect 2798 3819 2814 3853
rect 2614 3803 2814 3819
rect 2872 3853 3072 3900
rect 2872 3819 2888 3853
rect 3056 3819 3072 3853
rect 2872 3803 3072 3819
rect 3130 3853 3330 3900
rect 3130 3819 3146 3853
rect 3314 3819 3330 3853
rect 3130 3803 3330 3819
rect 3388 3853 3588 3900
rect 3388 3819 3404 3853
rect 3572 3819 3588 3853
rect 3388 3803 3588 3819
rect 3774 3853 3974 3900
rect 3774 3819 3790 3853
rect 3958 3819 3974 3853
rect 3774 3803 3974 3819
rect 414 3141 614 3157
rect 414 3107 430 3141
rect 598 3107 614 3141
rect 414 3060 614 3107
rect 794 3141 994 3157
rect 794 3107 810 3141
rect 978 3107 994 3141
rect 794 3060 994 3107
rect 1052 3141 1252 3157
rect 1052 3107 1068 3141
rect 1236 3107 1252 3141
rect 1052 3060 1252 3107
rect 1310 3141 1510 3157
rect 1310 3107 1326 3141
rect 1494 3107 1510 3141
rect 1310 3060 1510 3107
rect 1568 3141 1768 3157
rect 1568 3107 1584 3141
rect 1752 3107 1768 3141
rect 1568 3060 1768 3107
rect 1826 3141 2026 3157
rect 1826 3107 1842 3141
rect 2010 3107 2026 3141
rect 1826 3060 2026 3107
rect 2084 3141 2284 3157
rect 2084 3107 2100 3141
rect 2268 3107 2284 3141
rect 2084 3060 2284 3107
rect 2342 3141 2542 3157
rect 2342 3107 2358 3141
rect 2526 3107 2542 3141
rect 2342 3060 2542 3107
rect 2600 3141 2800 3157
rect 2600 3107 2616 3141
rect 2784 3107 2800 3141
rect 2600 3060 2800 3107
rect 2974 3141 3174 3157
rect 2974 3107 2990 3141
rect 3158 3107 3174 3141
rect 2974 3060 3174 3107
rect 414 2613 614 2660
rect 414 2579 430 2613
rect 598 2579 614 2613
rect 414 2563 614 2579
rect 794 2613 994 2660
rect 794 2579 810 2613
rect 978 2579 994 2613
rect 794 2563 994 2579
rect 1052 2613 1252 2660
rect 1052 2579 1068 2613
rect 1236 2579 1252 2613
rect 1052 2563 1252 2579
rect 1310 2613 1510 2660
rect 1310 2579 1326 2613
rect 1494 2579 1510 2613
rect 1310 2563 1510 2579
rect 1568 2613 1768 2660
rect 1568 2579 1584 2613
rect 1752 2579 1768 2613
rect 1568 2563 1768 2579
rect 1826 2613 2026 2660
rect 1826 2579 1842 2613
rect 2010 2579 2026 2613
rect 1826 2563 2026 2579
rect 2084 2613 2284 2660
rect 2084 2579 2100 2613
rect 2268 2579 2284 2613
rect 2084 2563 2284 2579
rect 2342 2613 2542 2660
rect 2342 2579 2358 2613
rect 2526 2579 2542 2613
rect 2342 2563 2542 2579
rect 2600 2613 2800 2660
rect 2600 2579 2616 2613
rect 2784 2579 2800 2613
rect 2600 2563 2800 2579
rect 2974 2613 3174 2660
rect 2974 2579 2990 2613
rect 3158 2579 3174 2613
rect 2974 2563 3174 2579
rect 5822 5363 6022 5379
rect 5822 5329 5838 5363
rect 6006 5329 6022 5363
rect 5822 5282 6022 5329
rect 6080 5363 6280 5379
rect 6080 5329 6096 5363
rect 6264 5329 6280 5363
rect 6080 5282 6280 5329
rect 6338 5363 6538 5379
rect 6338 5329 6354 5363
rect 6522 5329 6538 5363
rect 6338 5282 6538 5329
rect 6596 5363 6796 5379
rect 6596 5329 6612 5363
rect 6780 5329 6796 5363
rect 6596 5282 6796 5329
rect 6982 5363 7182 5379
rect 6982 5329 6998 5363
rect 7166 5329 7182 5363
rect 6982 5282 7182 5329
rect 7240 5363 7440 5379
rect 7240 5329 7256 5363
rect 7424 5329 7440 5363
rect 7240 5282 7440 5329
rect 7498 5363 7698 5379
rect 7498 5329 7514 5363
rect 7682 5329 7698 5363
rect 7498 5282 7698 5329
rect 7756 5363 7956 5379
rect 7756 5329 7772 5363
rect 7940 5329 7956 5363
rect 7756 5282 7956 5329
rect 8014 5363 8214 5379
rect 8014 5329 8030 5363
rect 8198 5329 8214 5363
rect 8014 5282 8214 5329
rect 8272 5363 8472 5379
rect 8272 5329 8288 5363
rect 8456 5329 8472 5363
rect 8272 5282 8472 5329
rect 8530 5363 8730 5379
rect 8530 5329 8546 5363
rect 8714 5329 8730 5363
rect 8530 5282 8730 5329
rect 8902 5363 9102 5379
rect 8902 5329 8918 5363
rect 9086 5329 9102 5363
rect 8902 5282 9102 5329
rect 9160 5363 9360 5379
rect 9160 5329 9176 5363
rect 9344 5329 9360 5363
rect 9160 5282 9360 5329
rect 9418 5363 9618 5379
rect 9418 5329 9434 5363
rect 9602 5329 9618 5363
rect 9418 5282 9618 5329
rect 9676 5363 9876 5379
rect 9676 5329 9692 5363
rect 9860 5329 9876 5363
rect 9676 5282 9876 5329
rect 9934 5363 10134 5379
rect 9934 5329 9950 5363
rect 10118 5329 10134 5363
rect 9934 5282 10134 5329
rect 10192 5363 10392 5379
rect 10192 5329 10208 5363
rect 10376 5329 10392 5363
rect 10192 5282 10392 5329
rect 10450 5363 10650 5379
rect 10450 5329 10466 5363
rect 10634 5329 10650 5363
rect 10450 5282 10650 5329
rect 10822 5363 11022 5379
rect 10822 5329 10838 5363
rect 11006 5329 11022 5363
rect 10822 5282 11022 5329
rect 11080 5363 11280 5379
rect 11080 5329 11096 5363
rect 11264 5329 11280 5363
rect 11080 5282 11280 5329
rect 11338 5363 11538 5379
rect 11338 5329 11354 5363
rect 11522 5329 11538 5363
rect 11338 5282 11538 5329
rect 11596 5363 11796 5379
rect 11596 5329 11612 5363
rect 11780 5329 11796 5363
rect 11596 5282 11796 5329
rect 6982 5035 7182 5082
rect 6982 5001 6998 5035
rect 7166 5001 7182 5035
rect 6982 4985 7182 5001
rect 7240 5035 7440 5082
rect 7240 5001 7256 5035
rect 7424 5001 7440 5035
rect 7240 4985 7440 5001
rect 7498 5035 7698 5082
rect 7498 5001 7514 5035
rect 7682 5001 7698 5035
rect 7498 4985 7698 5001
rect 7756 5035 7956 5082
rect 7756 5001 7772 5035
rect 7940 5001 7956 5035
rect 7756 4985 7956 5001
rect 8014 5035 8214 5082
rect 8014 5001 8030 5035
rect 8198 5001 8214 5035
rect 8014 4985 8214 5001
rect 8272 5035 8472 5082
rect 8272 5001 8288 5035
rect 8456 5001 8472 5035
rect 8272 4985 8472 5001
rect 8530 5035 8730 5082
rect 8530 5001 8546 5035
rect 8714 5001 8730 5035
rect 8530 4985 8730 5001
rect 8902 5035 9102 5082
rect 8902 5001 8918 5035
rect 9086 5001 9102 5035
rect 8902 4985 9102 5001
rect 9160 5035 9360 5082
rect 9160 5001 9176 5035
rect 9344 5001 9360 5035
rect 9160 4985 9360 5001
rect 9418 5035 9618 5082
rect 9418 5001 9434 5035
rect 9602 5001 9618 5035
rect 9418 4985 9618 5001
rect 9676 5035 9876 5082
rect 9676 5001 9692 5035
rect 9860 5001 9876 5035
rect 9676 4985 9876 5001
rect 9934 5035 10134 5082
rect 9934 5001 9950 5035
rect 10118 5001 10134 5035
rect 9934 4985 10134 5001
rect 10192 5035 10392 5082
rect 10192 5001 10208 5035
rect 10376 5001 10392 5035
rect 10192 4985 10392 5001
rect 10450 5035 10650 5082
rect 10450 5001 10466 5035
rect 10634 5001 10650 5035
rect 10450 4985 10650 5001
rect 5822 2235 6022 2282
rect 5822 2201 5838 2235
rect 6006 2201 6022 2235
rect 5822 2185 6022 2201
rect 6080 2235 6280 2282
rect 6080 2201 6096 2235
rect 6264 2201 6280 2235
rect 6080 2185 6280 2201
rect 6338 2235 6538 2282
rect 6338 2201 6354 2235
rect 6522 2201 6538 2235
rect 6338 2185 6538 2201
rect 6596 2235 6796 2282
rect 6596 2201 6612 2235
rect 6780 2201 6796 2235
rect 6596 2185 6796 2201
rect 8768 4682 8834 4698
rect 8768 4648 8784 4682
rect 8818 4648 8834 4682
rect 8690 4610 8720 4636
rect 8768 4632 8834 4648
rect 8960 4682 9026 4698
rect 8960 4648 8976 4682
rect 9010 4648 9026 4682
rect 8786 4610 8816 4632
rect 8882 4610 8912 4636
rect 8960 4632 9026 4648
rect 8978 4610 9008 4632
rect 8690 4288 8720 4310
rect 8672 4272 8738 4288
rect 8786 4284 8816 4310
rect 8882 4288 8912 4310
rect 8672 4238 8688 4272
rect 8722 4238 8738 4272
rect 8672 4222 8738 4238
rect 8864 4272 8930 4288
rect 8978 4284 9008 4310
rect 8864 4238 8880 4272
rect 8914 4238 8930 4272
rect 8864 4222 8930 4238
rect 7666 3962 7866 3978
rect 7666 3928 7682 3962
rect 7850 3928 7866 3962
rect 7666 3890 7866 3928
rect 7924 3962 8124 3978
rect 7924 3928 7940 3962
rect 8108 3928 8124 3962
rect 7924 3890 8124 3928
rect 8182 3962 8382 3978
rect 8182 3928 8198 3962
rect 8366 3928 8382 3962
rect 8182 3890 8382 3928
rect 8440 3962 8640 3978
rect 8440 3928 8456 3962
rect 8624 3928 8640 3962
rect 8440 3890 8640 3928
rect 8826 3902 9026 3918
rect 8826 3868 8842 3902
rect 9010 3868 9026 3902
rect 8826 3830 9026 3868
rect 9084 3902 9284 3918
rect 9084 3868 9100 3902
rect 9268 3868 9284 3902
rect 9084 3830 9284 3868
rect 9342 3902 9542 3918
rect 9342 3868 9358 3902
rect 9526 3868 9542 3902
rect 9342 3830 9542 3868
rect 9600 3902 9800 3918
rect 9600 3868 9616 3902
rect 9784 3868 9800 3902
rect 9600 3830 9800 3868
rect 9858 3902 10058 3918
rect 9858 3868 9874 3902
rect 10042 3868 10058 3902
rect 9858 3830 10058 3868
rect 10116 3902 10316 3918
rect 10116 3868 10132 3902
rect 10300 3868 10316 3902
rect 10116 3830 10316 3868
rect 7666 3652 7866 3690
rect 7666 3618 7682 3652
rect 7850 3618 7866 3652
rect 7666 3602 7866 3618
rect 7924 3652 8124 3690
rect 7924 3618 7940 3652
rect 8108 3618 8124 3652
rect 7924 3602 8124 3618
rect 8182 3652 8382 3690
rect 8182 3618 8198 3652
rect 8366 3618 8382 3652
rect 8182 3602 8382 3618
rect 8440 3652 8640 3690
rect 8440 3618 8456 3652
rect 8624 3618 8640 3652
rect 8440 3602 8640 3618
rect 8826 2792 9026 2830
rect 8826 2758 8842 2792
rect 9010 2758 9026 2792
rect 8826 2742 9026 2758
rect 9084 2792 9284 2830
rect 9084 2758 9100 2792
rect 9268 2758 9284 2792
rect 9084 2742 9284 2758
rect 9342 2792 9542 2830
rect 9342 2758 9358 2792
rect 9526 2758 9542 2792
rect 9342 2742 9542 2758
rect 9600 2792 9800 2830
rect 9600 2758 9616 2792
rect 9784 2758 9800 2792
rect 9600 2742 9800 2758
rect 9858 2792 10058 2830
rect 9858 2758 9874 2792
rect 10042 2758 10058 2792
rect 9858 2742 10058 2758
rect 10116 2792 10316 2830
rect 10116 2758 10132 2792
rect 10300 2758 10316 2792
rect 10116 2742 10316 2758
rect 10822 2235 11022 2282
rect 10822 2201 10838 2235
rect 11006 2201 11022 2235
rect 10822 2185 11022 2201
rect 11080 2235 11280 2282
rect 11080 2201 11096 2235
rect 11264 2201 11280 2235
rect 11080 2185 11280 2201
rect 11338 2235 11538 2282
rect 11338 2201 11354 2235
rect 11522 2201 11538 2235
rect 11338 2185 11538 2201
rect 11596 2235 11796 2282
rect 11596 2201 11612 2235
rect 11780 2201 11796 2235
rect 11596 2185 11796 2201
rect 218 1944 418 1960
rect 218 1910 234 1944
rect 402 1910 418 1944
rect 218 1872 418 1910
rect 598 1944 798 1960
rect 598 1910 614 1944
rect 782 1910 798 1944
rect 598 1872 798 1910
rect 978 1944 1178 1960
rect 978 1910 994 1944
rect 1162 1910 1178 1944
rect 978 1872 1178 1910
rect 1358 1944 1558 1960
rect 1358 1910 1374 1944
rect 1542 1910 1558 1944
rect 1358 1872 1558 1910
rect 1738 1944 1938 1960
rect 1738 1910 1754 1944
rect 1922 1910 1938 1944
rect 1738 1872 1938 1910
rect 2118 1944 2318 1960
rect 2118 1910 2134 1944
rect 2302 1910 2318 1944
rect 2118 1872 2318 1910
rect 2498 1944 2698 1960
rect 2498 1910 2514 1944
rect 2682 1910 2698 1944
rect 2498 1872 2698 1910
rect 2878 1944 3078 1960
rect 2878 1910 2894 1944
rect 3062 1910 3078 1944
rect 2878 1872 3078 1910
rect 218 1634 418 1672
rect 218 1600 234 1634
rect 402 1600 418 1634
rect 218 1584 418 1600
rect 598 1634 798 1672
rect 598 1600 614 1634
rect 782 1600 798 1634
rect 598 1584 798 1600
rect 978 1634 1178 1672
rect 978 1600 994 1634
rect 1162 1600 1178 1634
rect 978 1584 1178 1600
rect 1358 1634 1558 1672
rect 1358 1600 1374 1634
rect 1542 1600 1558 1634
rect 1358 1584 1558 1600
rect 1738 1634 1938 1672
rect 1738 1600 1754 1634
rect 1922 1600 1938 1634
rect 1738 1584 1938 1600
rect 2118 1634 2318 1672
rect 2118 1600 2134 1634
rect 2302 1600 2318 1634
rect 2118 1584 2318 1600
rect 2498 1634 2698 1672
rect 2498 1600 2514 1634
rect 2682 1600 2698 1634
rect 2498 1584 2698 1600
rect 2878 1634 3078 1672
rect 2878 1600 2894 1634
rect 3062 1600 3078 1634
rect 2878 1584 3078 1600
rect 218 1526 418 1542
rect 218 1492 234 1526
rect 402 1492 418 1526
rect 218 1454 418 1492
rect 598 1526 798 1542
rect 598 1492 614 1526
rect 782 1492 798 1526
rect 598 1454 798 1492
rect 978 1526 1178 1542
rect 978 1492 994 1526
rect 1162 1492 1178 1526
rect 978 1454 1178 1492
rect 1358 1526 1558 1542
rect 1358 1492 1374 1526
rect 1542 1492 1558 1526
rect 1358 1454 1558 1492
rect 1738 1526 1938 1542
rect 1738 1492 1754 1526
rect 1922 1492 1938 1526
rect 1738 1454 1938 1492
rect 2118 1526 2318 1542
rect 2118 1492 2134 1526
rect 2302 1492 2318 1526
rect 2118 1454 2318 1492
rect 2498 1526 2698 1542
rect 2498 1492 2514 1526
rect 2682 1492 2698 1526
rect 2498 1454 2698 1492
rect 2878 1526 3078 1542
rect 2878 1492 2894 1526
rect 3062 1492 3078 1526
rect 2878 1454 3078 1492
rect 218 1216 418 1254
rect 218 1182 234 1216
rect 402 1182 418 1216
rect 218 1166 418 1182
rect 598 1216 798 1254
rect 598 1182 614 1216
rect 782 1182 798 1216
rect 598 1166 798 1182
rect 978 1216 1178 1254
rect 978 1182 994 1216
rect 1162 1182 1178 1216
rect 978 1166 1178 1182
rect 1358 1216 1558 1254
rect 1358 1182 1374 1216
rect 1542 1182 1558 1216
rect 1358 1166 1558 1182
rect 1738 1216 1938 1254
rect 1738 1182 1754 1216
rect 1922 1182 1938 1216
rect 1738 1166 1938 1182
rect 2118 1216 2318 1254
rect 2118 1182 2134 1216
rect 2302 1182 2318 1216
rect 2118 1166 2318 1182
rect 2498 1216 2698 1254
rect 2498 1182 2514 1216
rect 2682 1182 2698 1216
rect 2498 1166 2698 1182
rect 2878 1216 3078 1254
rect 2878 1182 2894 1216
rect 3062 1182 3078 1216
rect 2878 1166 3078 1182
rect 218 1108 418 1124
rect 218 1074 234 1108
rect 402 1074 418 1108
rect 218 1036 418 1074
rect 598 1108 798 1124
rect 598 1074 614 1108
rect 782 1074 798 1108
rect 598 1036 798 1074
rect 978 1108 1178 1124
rect 978 1074 994 1108
rect 1162 1074 1178 1108
rect 978 1036 1178 1074
rect 1358 1108 1558 1124
rect 1358 1074 1374 1108
rect 1542 1074 1558 1108
rect 1358 1036 1558 1074
rect 1738 1108 1938 1124
rect 1738 1074 1754 1108
rect 1922 1074 1938 1108
rect 1738 1036 1938 1074
rect 2118 1108 2318 1124
rect 2118 1074 2134 1108
rect 2302 1074 2318 1108
rect 2118 1036 2318 1074
rect 2498 1108 2698 1124
rect 2498 1074 2514 1108
rect 2682 1074 2698 1108
rect 2498 1036 2698 1074
rect 2878 1108 3078 1124
rect 2878 1074 2894 1108
rect 3062 1074 3078 1108
rect 2878 1036 3078 1074
rect 218 798 418 836
rect 218 764 234 798
rect 402 764 418 798
rect 218 748 418 764
rect 598 798 798 836
rect 598 764 614 798
rect 782 764 798 798
rect 598 748 798 764
rect 978 798 1178 836
rect 978 764 994 798
rect 1162 764 1178 798
rect 978 748 1178 764
rect 1358 798 1558 836
rect 1358 764 1374 798
rect 1542 764 1558 798
rect 1358 748 1558 764
rect 1738 798 1938 836
rect 1738 764 1754 798
rect 1922 764 1938 798
rect 1738 748 1938 764
rect 2118 798 2318 836
rect 2118 764 2134 798
rect 2302 764 2318 798
rect 2118 748 2318 764
rect 2498 798 2698 836
rect 2498 764 2514 798
rect 2682 764 2698 798
rect 2498 748 2698 764
rect 2878 798 3078 836
rect 2878 764 2894 798
rect 3062 764 3078 798
rect 2878 748 3078 764
rect 218 690 418 706
rect 218 656 234 690
rect 402 656 418 690
rect 218 618 418 656
rect 598 690 798 706
rect 598 656 614 690
rect 782 656 798 690
rect 598 618 798 656
rect 978 690 1178 706
rect 978 656 994 690
rect 1162 656 1178 690
rect 978 618 1178 656
rect 1358 690 1558 706
rect 1358 656 1374 690
rect 1542 656 1558 690
rect 1358 618 1558 656
rect 1738 690 1938 706
rect 1738 656 1754 690
rect 1922 656 1938 690
rect 1738 618 1938 656
rect 2118 690 2318 706
rect 2118 656 2134 690
rect 2302 656 2318 690
rect 2118 618 2318 656
rect 2498 690 2698 706
rect 2498 656 2514 690
rect 2682 656 2698 690
rect 2498 618 2698 656
rect 2878 690 3078 706
rect 2878 656 2894 690
rect 3062 656 3078 690
rect 2878 618 3078 656
rect 218 380 418 418
rect 218 346 234 380
rect 402 346 418 380
rect 218 330 418 346
rect 598 380 798 418
rect 598 346 614 380
rect 782 346 798 380
rect 598 330 798 346
rect 978 380 1178 418
rect 978 346 994 380
rect 1162 346 1178 380
rect 978 330 1178 346
rect 1358 380 1558 418
rect 1358 346 1374 380
rect 1542 346 1558 380
rect 1358 330 1558 346
rect 1738 380 1938 418
rect 1738 346 1754 380
rect 1922 346 1938 380
rect 1738 330 1938 346
rect 2118 380 2318 418
rect 2118 346 2134 380
rect 2302 346 2318 380
rect 2118 330 2318 346
rect 2498 380 2698 418
rect 2498 346 2514 380
rect 2682 346 2698 380
rect 2498 330 2698 346
rect 2878 380 3078 418
rect 2878 346 2894 380
rect 3062 346 3078 380
rect 2878 330 3078 346
rect 14677 1299 14707 1325
rect 14761 1299 14791 1325
rect 15028 1305 15058 1331
rect 15120 1305 15150 1331
rect 15219 1305 15249 1331
rect 15359 1305 15389 1331
rect 15456 1305 15486 1331
rect 15653 1305 15683 1331
rect 15752 1305 15782 1331
rect 15838 1305 15868 1331
rect 15922 1305 15952 1331
rect 16030 1305 16060 1331
rect 16114 1305 16144 1331
rect 16278 1305 16308 1331
rect 16497 1305 16527 1331
rect 16594 1305 16624 1331
rect 14677 1156 14707 1171
rect 14644 1126 14707 1156
rect 14644 1073 14674 1126
rect 14761 1082 14791 1171
rect 15028 1134 15058 1221
rect 15120 1183 15150 1221
rect 14620 1057 14674 1073
rect 14620 1023 14630 1057
rect 14664 1023 14674 1057
rect 14716 1072 14791 1082
rect 14716 1038 14732 1072
rect 14766 1038 14791 1072
rect 14929 1118 15058 1134
rect 15104 1173 15170 1183
rect 15104 1139 15120 1173
rect 15154 1139 15170 1173
rect 15104 1129 15170 1139
rect 14929 1084 14939 1118
rect 14973 1104 15058 1118
rect 14973 1084 15046 1104
rect 15219 1087 15249 1221
rect 15359 1163 15389 1221
rect 15359 1147 15414 1163
rect 15359 1113 15369 1147
rect 15403 1113 15414 1147
rect 15359 1097 15414 1113
rect 14929 1068 15046 1084
rect 14716 1028 14791 1038
rect 14620 1007 14674 1023
rect 14644 984 14674 1007
rect 14644 954 14707 984
rect 14677 939 14707 954
rect 14761 939 14791 1028
rect 15016 939 15046 1068
rect 15111 1057 15249 1087
rect 15111 1027 15142 1057
rect 15088 1011 15142 1027
rect 15088 977 15098 1011
rect 15132 977 15142 1011
rect 15088 961 15142 977
rect 15184 1005 15250 1015
rect 15184 971 15200 1005
rect 15234 971 15250 1005
rect 15184 961 15250 971
rect 15111 927 15141 961
rect 15207 927 15237 961
rect 15373 939 15403 1097
rect 15456 1027 15486 1221
rect 15653 1122 15683 1137
rect 15577 1092 15683 1122
rect 15577 1075 15607 1092
rect 15541 1059 15607 1075
rect 15445 1011 15499 1027
rect 15445 977 15455 1011
rect 15489 977 15499 1011
rect 15541 1025 15551 1059
rect 15585 1025 15607 1059
rect 15752 1087 15782 1221
rect 15838 1189 15868 1221
rect 15824 1173 15878 1189
rect 15824 1139 15834 1173
rect 15868 1139 15878 1173
rect 15824 1123 15878 1139
rect 15752 1075 15802 1087
rect 15752 1063 15815 1075
rect 15752 1057 15839 1063
rect 15773 1047 15839 1057
rect 15773 1045 15795 1047
rect 15541 1009 15607 1025
rect 15577 983 15607 1009
rect 15676 999 15743 1015
rect 15445 961 15499 977
rect 15445 939 15475 961
rect 15676 965 15699 999
rect 15733 965 15743 999
rect 15676 949 15743 965
rect 15785 1013 15795 1045
rect 15829 1013 15839 1047
rect 15785 997 15839 1013
rect 15922 1037 15952 1221
rect 16030 1065 16060 1221
rect 16114 1173 16144 1221
rect 16102 1157 16156 1173
rect 16102 1123 16112 1157
rect 16146 1123 16156 1157
rect 16102 1107 16156 1123
rect 16025 1049 16079 1065
rect 15922 1021 15983 1037
rect 15922 1001 15939 1021
rect 15676 927 15706 949
rect 15785 927 15815 997
rect 15881 987 15939 1001
rect 15973 987 15983 1021
rect 16025 1015 16035 1049
rect 16069 1015 16079 1049
rect 16025 999 16079 1015
rect 15881 971 15983 987
rect 15881 939 15911 971
rect 16030 939 16060 999
rect 16121 939 16151 1107
rect 16497 1141 16527 1177
rect 16486 1111 16527 1141
rect 16278 1073 16308 1105
rect 16486 1073 16516 1111
rect 16594 1073 16624 1105
rect 16207 1057 16516 1073
rect 16207 1023 16235 1057
rect 16269 1023 16516 1057
rect 16207 1007 16516 1023
rect 16565 1057 16624 1073
rect 16565 1023 16575 1057
rect 16609 1023 16624 1057
rect 16565 1007 16624 1023
rect 16309 985 16339 1007
rect 16486 984 16516 1007
rect 16594 985 16624 1007
rect 17192 1834 17258 1850
rect 17192 1800 17208 1834
rect 17242 1800 17258 1834
rect 17192 1784 17258 1800
rect 17210 1753 17240 1784
rect 17210 1122 17240 1153
rect 17192 1106 17258 1122
rect 17192 1072 17208 1106
rect 17242 1072 17258 1106
rect 17192 1056 17258 1072
rect 16486 954 16527 984
rect 16497 939 16527 954
rect 14677 829 14707 855
rect 14761 829 14791 855
rect 15016 829 15046 855
rect 15111 829 15141 855
rect 15207 829 15237 855
rect 15373 829 15403 855
rect 15445 829 15475 855
rect 15577 829 15607 855
rect 15676 829 15706 855
rect 15785 829 15815 855
rect 15881 829 15911 855
rect 16030 829 16060 855
rect 16121 829 16151 855
rect 16309 829 16339 855
rect 16497 829 16527 855
rect 16594 829 16624 855
rect 17192 746 17258 762
rect 17192 712 17208 746
rect 17242 712 17258 746
rect 17192 696 17258 712
rect 17210 674 17240 696
rect 17210 452 17240 474
rect 17192 436 17258 452
rect 17192 402 17208 436
rect 17242 402 17258 436
rect 17192 386 17258 402
<< polycont >>
rect 1830 5027 1998 5061
rect 2210 5027 2378 5061
rect 2590 5027 3558 5061
rect 3770 5027 3938 5061
rect 1830 4499 1998 4533
rect 2210 4499 2378 4533
rect 2590 4499 3558 4533
rect 3770 4499 3938 4533
rect 450 4347 618 4381
rect 830 4347 998 4381
rect 1088 4347 1256 4381
rect 1470 4347 1638 4381
rect 1728 4347 1896 4381
rect 1986 4347 2154 4381
rect 2244 4347 2412 4381
rect 2630 4347 2798 4381
rect 2888 4347 3056 4381
rect 3146 4347 3314 4381
rect 3404 4347 3572 4381
rect 3790 4347 3958 4381
rect 450 3819 618 3853
rect 830 3819 998 3853
rect 1088 3819 1256 3853
rect 1470 3819 1638 3853
rect 1728 3819 1896 3853
rect 1986 3819 2154 3853
rect 2244 3819 2412 3853
rect 2630 3819 2798 3853
rect 2888 3819 3056 3853
rect 3146 3819 3314 3853
rect 3404 3819 3572 3853
rect 3790 3819 3958 3853
rect 430 3107 598 3141
rect 810 3107 978 3141
rect 1068 3107 1236 3141
rect 1326 3107 1494 3141
rect 1584 3107 1752 3141
rect 1842 3107 2010 3141
rect 2100 3107 2268 3141
rect 2358 3107 2526 3141
rect 2616 3107 2784 3141
rect 2990 3107 3158 3141
rect 430 2579 598 2613
rect 810 2579 978 2613
rect 1068 2579 1236 2613
rect 1326 2579 1494 2613
rect 1584 2579 1752 2613
rect 1842 2579 2010 2613
rect 2100 2579 2268 2613
rect 2358 2579 2526 2613
rect 2616 2579 2784 2613
rect 2990 2579 3158 2613
rect 5838 5329 6006 5363
rect 6096 5329 6264 5363
rect 6354 5329 6522 5363
rect 6612 5329 6780 5363
rect 6998 5329 7166 5363
rect 7256 5329 7424 5363
rect 7514 5329 7682 5363
rect 7772 5329 7940 5363
rect 8030 5329 8198 5363
rect 8288 5329 8456 5363
rect 8546 5329 8714 5363
rect 8918 5329 9086 5363
rect 9176 5329 9344 5363
rect 9434 5329 9602 5363
rect 9692 5329 9860 5363
rect 9950 5329 10118 5363
rect 10208 5329 10376 5363
rect 10466 5329 10634 5363
rect 10838 5329 11006 5363
rect 11096 5329 11264 5363
rect 11354 5329 11522 5363
rect 11612 5329 11780 5363
rect 6998 5001 7166 5035
rect 7256 5001 7424 5035
rect 7514 5001 7682 5035
rect 7772 5001 7940 5035
rect 8030 5001 8198 5035
rect 8288 5001 8456 5035
rect 8546 5001 8714 5035
rect 8918 5001 9086 5035
rect 9176 5001 9344 5035
rect 9434 5001 9602 5035
rect 9692 5001 9860 5035
rect 9950 5001 10118 5035
rect 10208 5001 10376 5035
rect 10466 5001 10634 5035
rect 5838 2201 6006 2235
rect 6096 2201 6264 2235
rect 6354 2201 6522 2235
rect 6612 2201 6780 2235
rect 8784 4648 8818 4682
rect 8976 4648 9010 4682
rect 8688 4238 8722 4272
rect 8880 4238 8914 4272
rect 7682 3928 7850 3962
rect 7940 3928 8108 3962
rect 8198 3928 8366 3962
rect 8456 3928 8624 3962
rect 8842 3868 9010 3902
rect 9100 3868 9268 3902
rect 9358 3868 9526 3902
rect 9616 3868 9784 3902
rect 9874 3868 10042 3902
rect 10132 3868 10300 3902
rect 7682 3618 7850 3652
rect 7940 3618 8108 3652
rect 8198 3618 8366 3652
rect 8456 3618 8624 3652
rect 8842 2758 9010 2792
rect 9100 2758 9268 2792
rect 9358 2758 9526 2792
rect 9616 2758 9784 2792
rect 9874 2758 10042 2792
rect 10132 2758 10300 2792
rect 10838 2201 11006 2235
rect 11096 2201 11264 2235
rect 11354 2201 11522 2235
rect 11612 2201 11780 2235
rect 234 1910 402 1944
rect 614 1910 782 1944
rect 994 1910 1162 1944
rect 1374 1910 1542 1944
rect 1754 1910 1922 1944
rect 2134 1910 2302 1944
rect 2514 1910 2682 1944
rect 2894 1910 3062 1944
rect 234 1600 402 1634
rect 614 1600 782 1634
rect 994 1600 1162 1634
rect 1374 1600 1542 1634
rect 1754 1600 1922 1634
rect 2134 1600 2302 1634
rect 2514 1600 2682 1634
rect 2894 1600 3062 1634
rect 234 1492 402 1526
rect 614 1492 782 1526
rect 994 1492 1162 1526
rect 1374 1492 1542 1526
rect 1754 1492 1922 1526
rect 2134 1492 2302 1526
rect 2514 1492 2682 1526
rect 2894 1492 3062 1526
rect 234 1182 402 1216
rect 614 1182 782 1216
rect 994 1182 1162 1216
rect 1374 1182 1542 1216
rect 1754 1182 1922 1216
rect 2134 1182 2302 1216
rect 2514 1182 2682 1216
rect 2894 1182 3062 1216
rect 234 1074 402 1108
rect 614 1074 782 1108
rect 994 1074 1162 1108
rect 1374 1074 1542 1108
rect 1754 1074 1922 1108
rect 2134 1074 2302 1108
rect 2514 1074 2682 1108
rect 2894 1074 3062 1108
rect 234 764 402 798
rect 614 764 782 798
rect 994 764 1162 798
rect 1374 764 1542 798
rect 1754 764 1922 798
rect 2134 764 2302 798
rect 2514 764 2682 798
rect 2894 764 3062 798
rect 234 656 402 690
rect 614 656 782 690
rect 994 656 1162 690
rect 1374 656 1542 690
rect 1754 656 1922 690
rect 2134 656 2302 690
rect 2514 656 2682 690
rect 2894 656 3062 690
rect 234 346 402 380
rect 614 346 782 380
rect 994 346 1162 380
rect 1374 346 1542 380
rect 1754 346 1922 380
rect 2134 346 2302 380
rect 2514 346 2682 380
rect 2894 346 3062 380
rect 14630 1023 14664 1057
rect 14732 1038 14766 1072
rect 15120 1139 15154 1173
rect 14939 1084 14973 1118
rect 15369 1113 15403 1147
rect 15098 977 15132 1011
rect 15200 971 15234 1005
rect 15455 977 15489 1011
rect 15551 1025 15585 1059
rect 15834 1139 15868 1173
rect 15699 965 15733 999
rect 15795 1013 15829 1047
rect 16112 1123 16146 1157
rect 15939 987 15973 1021
rect 16035 1015 16069 1049
rect 16235 1023 16269 1057
rect 16575 1023 16609 1057
rect 17208 1800 17242 1834
rect 17208 1072 17242 1106
rect 17208 712 17242 746
rect 17208 402 17242 436
<< xpolycontact >>
rect 14550 5320 14620 5752
rect 14550 3988 14620 4420
rect 14716 5320 14786 5752
rect 14716 3988 14786 4420
rect 14882 5320 14952 5752
rect 14882 3988 14952 4420
rect 15048 5320 15118 5752
rect 15048 3988 15118 4420
rect 15214 5320 15284 5752
rect 15214 3988 15284 4420
rect 15380 5320 15450 5752
rect 15380 3988 15450 4420
rect 15546 5320 15616 5752
rect 15546 3988 15616 4420
rect 15712 5320 15782 5752
rect 15712 3988 15782 4420
rect 16024 5320 16094 5752
rect 16024 3988 16094 4420
rect 16190 5320 16260 5752
rect 16190 3988 16260 4420
rect 16356 5320 16426 5752
rect 16356 3988 16426 4420
rect 16522 5320 16592 5752
rect 16522 3988 16592 4420
rect 16688 5320 16758 5752
rect 16688 3988 16758 4420
rect 16854 5320 16924 5752
rect 16854 3988 16924 4420
rect 17020 5320 17090 5752
rect 17020 3988 17090 4420
rect 17186 5320 17256 5752
rect 17186 3988 17256 4420
rect 14600 3152 14670 3584
rect 14600 2320 14670 2752
rect 14766 3152 14836 3584
rect 14766 2320 14836 2752
rect 14932 3152 15002 3584
rect 14932 2320 15002 2752
rect 15098 3152 15168 3584
rect 15098 2320 15168 2752
rect 15264 3152 15334 3584
rect 15264 2320 15334 2752
rect 15430 3152 15500 3584
rect 15430 2320 15500 2752
rect 15596 3152 15666 3584
rect 15596 2320 15666 2752
rect 15762 3152 15832 3584
rect 15762 2320 15832 2752
<< xpolyres >>
rect 14550 4420 14620 5320
rect 14716 4420 14786 5320
rect 14882 4420 14952 5320
rect 15048 4420 15118 5320
rect 15214 4420 15284 5320
rect 15380 4420 15450 5320
rect 15546 4420 15616 5320
rect 15712 4420 15782 5320
rect 16024 4420 16094 5320
rect 16190 4420 16260 5320
rect 16356 4420 16426 5320
rect 16522 4420 16592 5320
rect 16688 4420 16758 5320
rect 16854 4420 16924 5320
rect 17020 4420 17090 5320
rect 17186 4420 17256 5320
rect 14600 2752 14670 3152
rect 14766 2752 14836 3152
rect 14932 2752 15002 3152
rect 15098 2752 15168 3152
rect 15264 2752 15334 3152
rect 15430 2752 15500 3152
rect 15596 2752 15666 3152
rect 15762 2752 15832 3152
<< locali >>
rect 14396 5870 14492 5904
rect 17420 5870 17516 5904
rect 14396 5808 14430 5870
rect 11848 5499 11948 5502
rect 5671 5465 5731 5499
rect 11885 5465 11948 5499
rect 5671 5439 5705 5465
rect 7071 5462 7105 5465
rect 10571 5462 10605 5465
rect 11848 5462 11948 5465
rect 243 5223 303 5257
rect 4137 5223 4197 5257
rect 243 5197 277 5223
rect 4163 5197 4197 5223
rect 1814 5027 1830 5061
rect 1998 5027 2014 5061
rect 2194 5027 2210 5061
rect 2378 5027 2394 5061
rect 2574 5027 2590 5061
rect 3558 5027 3574 5061
rect 3754 5027 3770 5061
rect 3938 5027 3954 5061
rect 1768 4968 1802 4984
rect 1768 4576 1802 4592
rect 2026 4968 2060 4984
rect 2026 4576 2060 4592
rect 2148 4968 2182 4984
rect 2148 4576 2182 4592
rect 2406 4968 2440 4984
rect 2406 4576 2440 4592
rect 2528 4968 2562 4984
rect 2528 4576 2562 4592
rect 3586 4968 3620 4984
rect 3586 4576 3620 4592
rect 3708 4968 3742 4984
rect 3708 4576 3742 4592
rect 3966 4968 4000 4984
rect 3966 4576 4000 4592
rect 1814 4499 1830 4533
rect 1998 4499 2014 4533
rect 2194 4499 2210 4533
rect 2378 4499 2394 4533
rect 2574 4499 2590 4533
rect 3558 4499 3574 4533
rect 3754 4499 3770 4533
rect 3938 4499 3954 4533
rect 434 4347 450 4381
rect 618 4347 634 4381
rect 814 4347 830 4381
rect 998 4347 1014 4381
rect 1072 4347 1088 4381
rect 1256 4347 1272 4381
rect 1454 4347 1470 4381
rect 1638 4347 1654 4381
rect 1712 4347 1728 4381
rect 1896 4347 1912 4381
rect 1970 4347 1986 4381
rect 2154 4347 2170 4381
rect 2228 4347 2244 4381
rect 2412 4347 2428 4381
rect 2614 4347 2630 4381
rect 2798 4347 2814 4381
rect 2872 4347 2888 4381
rect 3056 4347 3072 4381
rect 3130 4347 3146 4381
rect 3314 4347 3330 4381
rect 3388 4347 3404 4381
rect 3572 4347 3588 4381
rect 3774 4347 3790 4381
rect 3958 4347 3974 4381
rect 388 4288 422 4304
rect 388 3896 422 3912
rect 646 4288 680 4304
rect 646 3896 680 3912
rect 768 4288 802 4304
rect 768 3896 802 3912
rect 1026 4288 1060 4304
rect 1026 3896 1060 3912
rect 1284 4288 1318 4304
rect 1284 3896 1318 3912
rect 1408 4288 1442 4304
rect 1408 3896 1442 3912
rect 1666 4288 1700 4304
rect 1666 3896 1700 3912
rect 1924 4288 1958 4304
rect 1924 3896 1958 3912
rect 2182 4288 2216 4304
rect 2182 3896 2216 3912
rect 2440 4288 2474 4304
rect 2440 3896 2474 3912
rect 2568 4288 2602 4304
rect 2568 3896 2602 3912
rect 2826 4288 2860 4304
rect 2826 3896 2860 3912
rect 3084 4288 3118 4304
rect 3084 3896 3118 3912
rect 3342 4288 3376 4304
rect 3342 3896 3376 3912
rect 3600 4288 3634 4304
rect 3600 3896 3634 3912
rect 3728 4288 3762 4304
rect 3728 3896 3762 3912
rect 3986 4288 4020 4304
rect 3986 3896 4020 3912
rect 434 3819 450 3853
rect 618 3819 634 3853
rect 814 3819 830 3853
rect 998 3819 1014 3853
rect 1072 3819 1088 3853
rect 1256 3819 1272 3853
rect 1454 3819 1470 3853
rect 1638 3819 1654 3853
rect 1712 3819 1728 3853
rect 1896 3819 1912 3853
rect 1970 3819 1986 3853
rect 2154 3819 2170 3853
rect 2228 3819 2244 3853
rect 2412 3819 2428 3853
rect 2614 3819 2630 3853
rect 2798 3819 2814 3853
rect 2872 3819 2888 3853
rect 3056 3819 3072 3853
rect 3130 3819 3146 3853
rect 3314 3819 3330 3853
rect 3388 3819 3404 3853
rect 3572 3819 3588 3853
rect 3774 3819 3790 3853
rect 3958 3819 3974 3853
rect 243 3697 277 3723
rect 4163 3697 4197 3723
rect 243 3663 303 3697
rect 4137 3663 4197 3697
rect 203 3303 263 3337
rect 3297 3303 3357 3337
rect 203 3277 237 3303
rect 3323 3277 3357 3303
rect 414 3107 430 3141
rect 598 3107 614 3141
rect 794 3107 810 3141
rect 978 3107 994 3141
rect 1052 3107 1068 3141
rect 1236 3107 1252 3141
rect 1310 3107 1326 3141
rect 1494 3107 1510 3141
rect 1568 3107 1584 3141
rect 1752 3107 1768 3141
rect 1826 3107 1842 3141
rect 2010 3107 2026 3141
rect 2084 3107 2100 3141
rect 2268 3107 2284 3141
rect 2342 3107 2358 3141
rect 2526 3107 2542 3141
rect 2600 3107 2616 3141
rect 2784 3107 2800 3141
rect 2974 3107 2990 3141
rect 3158 3107 3174 3141
rect 368 3048 402 3064
rect 368 2656 402 2672
rect 626 3048 660 3064
rect 626 2656 660 2672
rect 748 3048 782 3064
rect 748 2656 782 2672
rect 1006 3048 1040 3064
rect 1006 2656 1040 2672
rect 1264 3048 1298 3064
rect 1264 2656 1298 2672
rect 1522 3048 1556 3064
rect 1522 2656 1556 2672
rect 1780 3048 1814 3064
rect 1780 2656 1814 2672
rect 2038 3048 2072 3064
rect 2038 2656 2072 2672
rect 2296 3048 2330 3064
rect 2296 2656 2330 2672
rect 2554 3048 2588 3064
rect 2554 2656 2588 2672
rect 2812 3048 2846 3064
rect 2812 2656 2846 2672
rect 2928 3048 2962 3064
rect 2928 2656 2962 2672
rect 3186 3048 3220 3064
rect 3186 2656 3220 2672
rect 414 2579 430 2613
rect 598 2579 614 2613
rect 794 2579 810 2613
rect 978 2579 994 2613
rect 1052 2579 1068 2613
rect 1236 2579 1252 2613
rect 1310 2579 1326 2613
rect 1494 2579 1510 2613
rect 1568 2579 1584 2613
rect 1752 2579 1768 2613
rect 1826 2579 1842 2613
rect 2010 2579 2026 2613
rect 2084 2579 2100 2613
rect 2268 2579 2284 2613
rect 2342 2579 2358 2613
rect 2526 2579 2542 2613
rect 2600 2579 2616 2613
rect 2784 2579 2800 2613
rect 2974 2579 2990 2613
rect 3158 2579 3174 2613
rect 203 2377 237 2403
rect 3323 2377 3357 2403
rect 203 2343 263 2377
rect 3297 2343 3357 2377
rect 11911 5439 11945 5462
rect 5822 5329 5838 5363
rect 6006 5329 6022 5363
rect 6080 5329 6096 5363
rect 6264 5329 6280 5363
rect 6338 5329 6354 5363
rect 6522 5329 6538 5363
rect 6596 5329 6612 5363
rect 6780 5329 6796 5363
rect 6982 5329 6998 5363
rect 7166 5329 7182 5363
rect 7240 5329 7256 5363
rect 7424 5329 7440 5363
rect 7498 5329 7514 5363
rect 7682 5329 7698 5363
rect 7756 5329 7772 5363
rect 7940 5329 7956 5363
rect 8014 5329 8030 5363
rect 8198 5329 8214 5363
rect 8272 5329 8288 5363
rect 8456 5329 8472 5363
rect 8530 5329 8546 5363
rect 8714 5329 8730 5363
rect 8902 5329 8918 5363
rect 9086 5329 9102 5363
rect 9160 5329 9176 5363
rect 9344 5329 9360 5363
rect 9418 5329 9434 5363
rect 9602 5329 9618 5363
rect 9676 5329 9692 5363
rect 9860 5329 9876 5363
rect 9934 5329 9950 5363
rect 10118 5329 10134 5363
rect 10192 5329 10208 5363
rect 10376 5329 10392 5363
rect 10450 5329 10466 5363
rect 10634 5329 10650 5363
rect 10822 5329 10838 5363
rect 11006 5329 11022 5363
rect 11080 5329 11096 5363
rect 11264 5329 11280 5363
rect 11338 5329 11354 5363
rect 11522 5329 11538 5363
rect 11596 5329 11612 5363
rect 11780 5329 11796 5363
rect 5776 5270 5810 5286
rect 5705 4845 5708 4879
rect 5776 2278 5810 2294
rect 6034 5270 6068 5286
rect 6034 2278 6068 2294
rect 6292 5270 6326 5286
rect 6292 2278 6326 2294
rect 6550 5270 6584 5286
rect 6550 2278 6584 2294
rect 6808 5270 6842 5286
rect 6936 5270 6970 5286
rect 6936 5078 6970 5094
rect 7194 5270 7228 5286
rect 7194 5078 7228 5094
rect 7452 5270 7486 5286
rect 7452 5078 7486 5094
rect 7710 5270 7744 5286
rect 7710 5078 7744 5094
rect 7968 5270 8002 5286
rect 7968 5078 8002 5094
rect 8226 5270 8260 5286
rect 8226 5078 8260 5094
rect 8484 5270 8518 5286
rect 8484 5078 8518 5094
rect 8742 5270 8776 5286
rect 8742 5078 8776 5094
rect 8856 5270 8890 5286
rect 8856 5078 8890 5094
rect 9114 5270 9148 5286
rect 9114 5078 9148 5094
rect 9372 5270 9406 5286
rect 9372 5078 9406 5094
rect 9630 5270 9664 5286
rect 9630 5078 9664 5094
rect 9888 5270 9922 5286
rect 9888 5078 9922 5094
rect 10146 5270 10180 5286
rect 10146 5078 10180 5094
rect 10404 5270 10438 5286
rect 10404 5078 10438 5094
rect 10662 5270 10696 5286
rect 10662 5078 10696 5094
rect 10776 5270 10810 5286
rect 6982 5001 6998 5035
rect 7166 5001 7182 5035
rect 7240 5001 7256 5035
rect 7424 5001 7440 5035
rect 7498 5001 7514 5035
rect 7682 5001 7698 5035
rect 7756 5001 7772 5035
rect 7940 5001 7956 5035
rect 8014 5001 8030 5035
rect 8198 5001 8214 5035
rect 8272 5001 8288 5035
rect 8456 5001 8472 5035
rect 8530 5001 8546 5035
rect 8714 5001 8730 5035
rect 8902 5001 8918 5035
rect 9160 5001 9176 5035
rect 9418 5001 9434 5035
rect 9676 5001 9692 5035
rect 9934 5001 9950 5035
rect 10192 5001 10208 5035
rect 10376 5001 10392 5035
rect 10450 5001 10466 5035
rect 6948 4879 7208 4882
rect 10671 4879 10705 4882
rect 6928 4845 7148 4879
rect 10528 4845 10705 4879
rect 6928 4842 7208 4845
rect 6928 4765 6965 4842
rect 10671 4802 10705 4845
rect 6808 2278 6842 2294
rect 6931 4762 6965 4765
rect 5822 2201 5838 2235
rect 6006 2201 6022 2235
rect 6080 2201 6096 2235
rect 6264 2201 6280 2235
rect 6338 2201 6354 2235
rect 6522 2201 6538 2235
rect 6596 2201 6612 2235
rect 6780 2201 6796 2235
rect 5671 2119 5705 2145
rect 7344 4732 7440 4766
rect 10368 4732 10464 4766
rect 7344 4670 7378 4732
rect 8768 4648 8784 4682
rect 8818 4648 8834 4682
rect 8960 4648 8976 4682
rect 9010 4648 9026 4682
rect 10430 4670 10464 4732
rect 8640 4598 8674 4614
rect 8640 4306 8674 4322
rect 8736 4598 8770 4614
rect 8736 4306 8770 4322
rect 8832 4598 8866 4614
rect 8832 4306 8866 4322
rect 8928 4598 8962 4614
rect 8928 4306 8962 4322
rect 9024 4598 9058 4614
rect 9024 4306 9058 4322
rect 8672 4238 8688 4272
rect 8722 4238 8738 4272
rect 8864 4238 8880 4272
rect 8914 4238 8930 4272
rect 7666 3928 7682 3962
rect 7850 3928 7866 3962
rect 7924 3928 7940 3962
rect 8108 3928 8124 3962
rect 8182 3928 8198 3962
rect 8366 3928 8382 3962
rect 8440 3928 8456 3962
rect 8624 3928 8640 3962
rect 7620 3878 7654 3894
rect 7620 3686 7654 3702
rect 7878 3878 7912 3894
rect 7878 3686 7912 3702
rect 8136 3878 8170 3894
rect 8136 3686 8170 3702
rect 8394 3878 8428 3894
rect 8394 3686 8428 3702
rect 8652 3878 8686 3894
rect 8826 3868 8842 3902
rect 9010 3868 9026 3902
rect 9084 3868 9100 3902
rect 9268 3868 9284 3902
rect 9342 3868 9358 3902
rect 9526 3868 9542 3902
rect 9600 3868 9616 3902
rect 9784 3868 9800 3902
rect 9858 3868 9874 3902
rect 10042 3868 10058 3902
rect 10116 3868 10132 3902
rect 10300 3868 10316 3902
rect 8652 3686 8686 3702
rect 8780 3818 8814 3834
rect 7666 3618 7682 3652
rect 7850 3618 7866 3652
rect 7924 3618 7940 3652
rect 8108 3618 8124 3652
rect 8182 3618 8198 3652
rect 8366 3618 8382 3652
rect 8440 3618 8456 3652
rect 8624 3618 8640 3652
rect 8780 2826 8814 2842
rect 9038 3818 9072 3834
rect 9038 2826 9072 2842
rect 9296 3818 9330 3834
rect 9296 2826 9330 2842
rect 9554 3818 9588 3834
rect 9554 2826 9588 2842
rect 9812 3818 9846 3834
rect 9812 2826 9846 2842
rect 10070 3818 10104 3834
rect 10070 2826 10104 2842
rect 10328 3818 10362 3834
rect 10328 2826 10362 2842
rect 8826 2758 8842 2792
rect 9010 2758 9026 2792
rect 9084 2758 9100 2792
rect 9268 2758 9284 2792
rect 9342 2758 9358 2792
rect 9526 2758 9542 2792
rect 9600 2758 9616 2792
rect 9784 2758 9800 2792
rect 9858 2758 9874 2792
rect 10042 2758 10058 2792
rect 10116 2758 10132 2792
rect 10300 2758 10316 2792
rect 7344 2652 7378 2714
rect 10430 2652 10464 2714
rect 7344 2618 7440 2652
rect 10368 2618 10464 2652
rect 6931 2119 6965 2145
rect 5671 2085 5731 2119
rect 6905 2085 6965 2119
rect 10776 2278 10810 2294
rect 11034 5270 11068 5286
rect 11034 2278 11068 2294
rect 11292 5270 11326 5286
rect 11292 2278 11326 2294
rect 11550 5270 11584 5286
rect 11550 2278 11584 2294
rect 11808 5270 11842 5286
rect 11908 4845 11911 4879
rect 11808 2278 11842 2294
rect 10822 2201 10838 2235
rect 11006 2201 11022 2235
rect 11080 2201 11096 2235
rect 11264 2201 11280 2235
rect 11338 2201 11354 2235
rect 11522 2201 11538 2235
rect 11596 2201 11612 2235
rect 11780 2201 11796 2235
rect 10671 2119 10705 2145
rect 17482 5808 17516 5870
rect 14396 2190 14430 2252
rect 16020 2190 16140 2200
rect 17482 2190 17516 2252
rect 14396 2156 14492 2190
rect 17420 2156 17516 2190
rect 11911 2119 11945 2145
rect 10671 2085 10731 2119
rect 11885 2085 11945 2119
rect 36 2010 132 2044
rect 3260 2010 3356 2044
rect 36 1948 70 2010
rect 3322 1948 3356 2010
rect 218 1910 234 1944
rect 402 1910 418 1944
rect 598 1910 614 1944
rect 782 1910 798 1944
rect 978 1910 994 1944
rect 1162 1910 1178 1944
rect 1358 1910 1374 1944
rect 1542 1910 1558 1944
rect 1738 1910 1754 1944
rect 1922 1910 1938 1944
rect 2118 1910 2134 1944
rect 2302 1910 2318 1944
rect 2498 1910 2514 1944
rect 2682 1910 2698 1944
rect 2878 1910 2894 1944
rect 3062 1910 3078 1944
rect 172 1860 206 1876
rect 172 1668 206 1684
rect 430 1860 464 1876
rect 430 1668 464 1684
rect 552 1860 586 1876
rect 552 1668 586 1684
rect 810 1860 844 1876
rect 810 1668 844 1684
rect 932 1860 966 1876
rect 932 1668 966 1684
rect 1190 1860 1224 1876
rect 1190 1668 1224 1684
rect 1312 1860 1346 1876
rect 1312 1668 1346 1684
rect 1570 1860 1604 1876
rect 1570 1668 1604 1684
rect 1692 1860 1726 1876
rect 1692 1668 1726 1684
rect 1950 1860 1984 1876
rect 1950 1668 1984 1684
rect 2072 1860 2106 1876
rect 2072 1668 2106 1684
rect 2330 1860 2364 1876
rect 2330 1668 2364 1684
rect 2452 1860 2486 1876
rect 2452 1668 2486 1684
rect 2710 1860 2744 1876
rect 2710 1668 2744 1684
rect 2832 1860 2866 1876
rect 2832 1668 2866 1684
rect 3090 1860 3124 1876
rect 3090 1668 3124 1684
rect 218 1600 234 1634
rect 402 1600 418 1634
rect 598 1600 614 1634
rect 782 1600 798 1634
rect 978 1600 994 1634
rect 1162 1600 1178 1634
rect 1358 1600 1374 1634
rect 1542 1600 1558 1634
rect 1738 1600 1754 1634
rect 1922 1600 1938 1634
rect 2118 1600 2134 1634
rect 2302 1600 2318 1634
rect 2498 1600 2514 1634
rect 2682 1600 2698 1634
rect 2878 1600 2894 1634
rect 3062 1600 3078 1634
rect 218 1492 234 1526
rect 402 1492 418 1526
rect 598 1492 614 1526
rect 782 1492 798 1526
rect 978 1492 994 1526
rect 1162 1492 1178 1526
rect 1358 1492 1374 1526
rect 1542 1492 1558 1526
rect 1738 1492 1754 1526
rect 1922 1492 1938 1526
rect 2118 1492 2134 1526
rect 2302 1492 2318 1526
rect 2498 1492 2514 1526
rect 2682 1492 2698 1526
rect 2878 1492 2894 1526
rect 3062 1492 3078 1526
rect 172 1442 206 1458
rect 172 1250 206 1266
rect 430 1442 464 1458
rect 430 1250 464 1266
rect 552 1442 586 1458
rect 552 1250 586 1266
rect 810 1442 844 1458
rect 810 1250 844 1266
rect 932 1442 966 1458
rect 932 1250 966 1266
rect 1190 1442 1224 1458
rect 1190 1250 1224 1266
rect 1312 1442 1346 1458
rect 1312 1250 1346 1266
rect 1570 1442 1604 1458
rect 1570 1250 1604 1266
rect 1692 1442 1726 1458
rect 1692 1250 1726 1266
rect 1950 1442 1984 1458
rect 1950 1250 1984 1266
rect 2072 1442 2106 1458
rect 2072 1250 2106 1266
rect 2330 1442 2364 1458
rect 2330 1250 2364 1266
rect 2452 1442 2486 1458
rect 2452 1250 2486 1266
rect 2710 1442 2744 1458
rect 2710 1250 2744 1266
rect 2832 1442 2866 1458
rect 2832 1250 2866 1266
rect 3090 1442 3124 1458
rect 3090 1250 3124 1266
rect 218 1182 234 1216
rect 402 1182 418 1216
rect 598 1182 614 1216
rect 782 1182 798 1216
rect 978 1182 994 1216
rect 1162 1182 1178 1216
rect 1358 1182 1374 1216
rect 1542 1182 1558 1216
rect 1738 1182 1754 1216
rect 1922 1182 1938 1216
rect 2118 1182 2134 1216
rect 2302 1182 2318 1216
rect 2498 1182 2514 1216
rect 2682 1182 2698 1216
rect 2878 1182 2894 1216
rect 3062 1182 3078 1216
rect 218 1074 234 1108
rect 402 1074 418 1108
rect 598 1074 614 1108
rect 782 1074 798 1108
rect 978 1074 994 1108
rect 1162 1074 1178 1108
rect 1358 1074 1374 1108
rect 1542 1074 1558 1108
rect 1738 1074 1754 1108
rect 1922 1074 1938 1108
rect 2118 1074 2134 1108
rect 2302 1074 2318 1108
rect 2498 1074 2514 1108
rect 2682 1074 2698 1108
rect 2878 1074 2894 1108
rect 3062 1074 3078 1108
rect 172 1024 206 1040
rect 172 832 206 848
rect 430 1024 464 1040
rect 430 832 464 848
rect 552 1024 586 1040
rect 552 832 586 848
rect 810 1024 844 1040
rect 810 832 844 848
rect 932 1024 966 1040
rect 932 832 966 848
rect 1190 1024 1224 1040
rect 1190 832 1224 848
rect 1312 1024 1346 1040
rect 1312 832 1346 848
rect 1570 1024 1604 1040
rect 1570 832 1604 848
rect 1692 1024 1726 1040
rect 1692 832 1726 848
rect 1950 1024 1984 1040
rect 1950 832 1984 848
rect 2072 1024 2106 1040
rect 2072 832 2106 848
rect 2330 1024 2364 1040
rect 2330 832 2364 848
rect 2452 1024 2486 1040
rect 2452 832 2486 848
rect 2710 1024 2744 1040
rect 2710 832 2744 848
rect 2832 1024 2866 1040
rect 2832 832 2866 848
rect 3090 1024 3124 1040
rect 3090 832 3124 848
rect 218 764 234 798
rect 402 764 418 798
rect 598 764 614 798
rect 782 764 798 798
rect 978 764 994 798
rect 1162 764 1178 798
rect 1358 764 1374 798
rect 1542 764 1558 798
rect 1738 764 1754 798
rect 1922 764 1938 798
rect 2118 764 2134 798
rect 2302 764 2318 798
rect 2498 764 2514 798
rect 2682 764 2698 798
rect 2878 764 2894 798
rect 3062 764 3078 798
rect 218 656 234 690
rect 402 656 418 690
rect 598 656 614 690
rect 782 656 798 690
rect 978 656 994 690
rect 1162 656 1178 690
rect 1358 656 1374 690
rect 1542 656 1558 690
rect 1738 656 1754 690
rect 1922 656 1938 690
rect 2118 656 2134 690
rect 2302 656 2318 690
rect 2498 656 2514 690
rect 2682 656 2698 690
rect 2878 656 2894 690
rect 3062 656 3078 690
rect 172 606 206 622
rect 172 414 206 430
rect 430 606 464 622
rect 430 414 464 430
rect 552 606 586 622
rect 552 414 586 430
rect 810 606 844 622
rect 810 414 844 430
rect 932 606 966 622
rect 932 414 966 430
rect 1190 606 1224 622
rect 1190 414 1224 430
rect 1312 606 1346 622
rect 1312 414 1346 430
rect 1570 606 1604 622
rect 1570 414 1604 430
rect 1692 606 1726 622
rect 1692 414 1726 430
rect 1950 606 1984 622
rect 1950 414 1984 430
rect 2072 606 2106 622
rect 2072 414 2106 430
rect 2330 606 2364 622
rect 2330 414 2364 430
rect 2452 606 2486 622
rect 2452 414 2486 430
rect 2710 606 2744 622
rect 2710 414 2744 430
rect 2832 606 2866 622
rect 2832 414 2866 430
rect 3090 606 3124 622
rect 3090 414 3124 430
rect 218 346 234 380
rect 402 346 418 380
rect 598 346 614 380
rect 782 346 798 380
rect 978 346 994 380
rect 1162 346 1178 380
rect 1358 346 1374 380
rect 1542 346 1558 380
rect 1738 346 1754 380
rect 1922 346 1938 380
rect 2118 346 2134 380
rect 2302 346 2318 380
rect 2498 346 2514 380
rect 2682 346 2698 380
rect 2878 346 2894 380
rect 3062 346 3078 380
rect 36 230 70 292
rect 17050 1902 17146 1936
rect 17304 1902 17400 1936
rect 17050 1840 17084 1902
rect 14598 1335 14627 1369
rect 14661 1335 14719 1369
rect 14753 1335 14811 1369
rect 14845 1335 14903 1369
rect 14937 1335 14995 1369
rect 15029 1335 15087 1369
rect 15121 1335 15179 1369
rect 15213 1335 15271 1369
rect 15305 1335 15363 1369
rect 15397 1335 15455 1369
rect 15489 1335 15547 1369
rect 15581 1335 15639 1369
rect 15673 1335 15731 1369
rect 15765 1335 15823 1369
rect 15857 1335 15915 1369
rect 15949 1335 16007 1369
rect 16041 1335 16099 1369
rect 16133 1335 16191 1369
rect 16225 1335 16283 1369
rect 16317 1335 16375 1369
rect 16409 1335 16467 1369
rect 16501 1335 16559 1369
rect 16593 1335 16651 1369
rect 16685 1335 16714 1369
rect 14420 1300 14520 1310
rect 14420 1250 14430 1300
rect 14500 1250 14520 1300
rect 14420 1220 14520 1250
rect 14616 1285 14667 1301
rect 14616 1251 14633 1285
rect 14616 1217 14667 1251
rect 14701 1269 14767 1335
rect 14701 1235 14717 1269
rect 14751 1235 14767 1269
rect 14801 1285 14835 1301
rect 14616 1183 14633 1217
rect 14801 1217 14835 1251
rect 14667 1183 14766 1201
rect 14616 1167 14766 1183
rect 14616 1080 14686 1133
rect 14616 1020 14620 1080
rect 14660 1057 14686 1080
rect 14664 1023 14686 1057
rect 14660 1020 14686 1023
rect 14616 1003 14686 1020
rect 14720 1072 14766 1167
rect 14720 1063 14732 1072
rect 14754 1029 14766 1038
rect 14720 969 14766 1029
rect 14616 935 14766 969
rect 14616 927 14667 935
rect 14616 893 14633 927
rect 14801 927 14835 1165
rect 14869 1141 14934 1298
rect 14968 1293 15018 1335
rect 14968 1259 14984 1293
rect 14968 1243 15018 1259
rect 15052 1285 15102 1301
rect 15052 1251 15068 1285
rect 15052 1235 15102 1251
rect 15145 1291 15281 1301
rect 15145 1257 15161 1291
rect 15195 1257 15281 1291
rect 15396 1283 15462 1335
rect 15589 1293 15663 1335
rect 15145 1235 15281 1257
rect 15052 1209 15086 1235
rect 15007 1175 15086 1209
rect 15120 1199 15213 1201
rect 14881 1118 14973 1141
rect 14881 1084 14939 1118
rect 14881 990 14973 1084
rect 14881 950 14900 990
rect 14960 950 14973 990
rect 14881 931 14973 950
rect 14616 877 14667 893
rect 14701 867 14717 901
rect 14751 867 14767 901
rect 15007 903 15041 1175
rect 15120 1173 15179 1199
rect 15154 1165 15179 1173
rect 15154 1139 15213 1165
rect 15120 1123 15213 1139
rect 15075 1063 15145 1085
rect 15075 1029 15087 1063
rect 15121 1029 15145 1063
rect 15075 1011 15145 1029
rect 15075 977 15098 1011
rect 15132 977 15145 1011
rect 15075 961 15145 977
rect 15179 1005 15213 1123
rect 15247 1079 15281 1235
rect 15315 1267 15349 1283
rect 15396 1249 15412 1283
rect 15446 1249 15462 1283
rect 15496 1267 15530 1283
rect 15315 1215 15349 1233
rect 15589 1259 15609 1293
rect 15643 1259 15663 1293
rect 15589 1243 15663 1259
rect 15697 1285 15731 1301
rect 15496 1215 15530 1233
rect 15315 1181 15530 1215
rect 15697 1209 15731 1251
rect 15778 1292 15952 1301
rect 15778 1258 15794 1292
rect 15828 1258 15952 1292
rect 15778 1233 15952 1258
rect 15986 1293 16036 1335
rect 16020 1259 16036 1293
rect 16140 1293 16284 1335
rect 15986 1243 16036 1259
rect 16070 1267 16104 1283
rect 15619 1175 15731 1209
rect 15619 1147 15653 1175
rect 15353 1113 15369 1147
rect 15403 1113 15653 1147
rect 15792 1165 15803 1199
rect 15837 1173 15884 1199
rect 15792 1141 15834 1165
rect 15247 1059 15585 1079
rect 15247 1045 15551 1059
rect 15179 971 15200 1005
rect 15234 971 15250 1005
rect 15179 961 15250 971
rect 15284 903 15318 1045
rect 15359 995 15455 1011
rect 15393 961 15431 995
rect 15489 977 15517 1011
rect 15551 1009 15585 1025
rect 15465 961 15517 977
rect 15619 975 15653 1113
rect 14801 877 14835 893
rect 14701 825 14767 867
rect 14907 863 14923 897
rect 14957 863 14973 897
rect 15007 869 15056 903
rect 15090 869 15106 903
rect 15147 869 15163 903
rect 15197 869 15318 903
rect 15493 901 15559 917
rect 14907 825 14973 863
rect 15493 867 15509 901
rect 15543 867 15559 901
rect 15493 825 15559 867
rect 15601 897 15653 975
rect 15691 1139 15834 1141
rect 15868 1139 15884 1173
rect 15918 1157 15952 1233
rect 16140 1259 16156 1293
rect 16190 1259 16234 1293
rect 16268 1259 16284 1293
rect 16318 1285 16399 1301
rect 16550 1293 16584 1335
rect 16070 1225 16104 1233
rect 16352 1251 16399 1285
rect 16070 1191 16230 1225
rect 15691 1107 15826 1139
rect 15918 1123 16112 1157
rect 16146 1123 16162 1157
rect 15691 999 15733 1107
rect 15918 1105 15952 1123
rect 15691 965 15699 999
rect 15691 949 15733 965
rect 15767 1063 15837 1073
rect 15767 1047 15803 1063
rect 15767 1013 15795 1047
rect 15829 1013 15837 1029
rect 15767 949 15837 1013
rect 15871 1071 15952 1105
rect 15871 915 15905 1071
rect 16019 1058 16127 1089
rect 16196 1073 16230 1191
rect 16318 1217 16399 1251
rect 16352 1183 16399 1217
rect 16318 1149 16399 1183
rect 16352 1115 16399 1149
rect 16318 1099 16399 1115
rect 16196 1067 16285 1073
rect 16053 1049 16127 1058
rect 15939 1021 15983 1037
rect 15973 987 15983 1021
rect 16019 1015 16035 1024
rect 16069 1015 16127 1049
rect 15939 981 15983 987
rect 16079 995 16127 1015
rect 15939 947 16045 981
rect 15715 901 15905 915
rect 15601 863 15621 897
rect 15655 863 15671 897
rect 15715 867 15731 901
rect 15765 867 15905 901
rect 15715 859 15905 867
rect 15939 897 15977 913
rect 15939 863 15943 897
rect 16011 901 16045 947
rect 16113 961 16127 995
rect 16079 935 16127 961
rect 16161 1057 16285 1067
rect 16161 1023 16235 1057
rect 16269 1023 16285 1057
rect 16161 1007 16285 1023
rect 16161 972 16226 1007
rect 16333 973 16399 1099
rect 16161 917 16225 972
rect 16011 883 16161 901
rect 16195 883 16225 917
rect 16011 867 16225 883
rect 16265 940 16299 962
rect 15939 825 15977 863
rect 16265 825 16299 906
rect 16333 960 16349 973
rect 16383 960 16399 973
rect 16437 1259 16453 1293
rect 16487 1259 16503 1293
rect 16437 1225 16503 1259
rect 16437 1191 16453 1225
rect 16487 1191 16503 1225
rect 16437 1073 16503 1191
rect 16550 1225 16584 1259
rect 16550 1157 16584 1191
rect 16550 1107 16584 1123
rect 16634 1257 16685 1273
rect 16668 1223 16685 1257
rect 16634 1189 16685 1223
rect 16668 1155 16685 1189
rect 16634 1097 16685 1155
rect 16437 1057 16609 1073
rect 16437 1023 16575 1057
rect 16437 1007 16609 1023
rect 16643 1060 16685 1097
rect 17366 1840 17400 1902
rect 17192 1800 17208 1834
rect 17242 1800 17258 1834
rect 17164 1741 17198 1757
rect 17164 1149 17198 1165
rect 17252 1741 17286 1757
rect 17252 1149 17286 1165
rect 17192 1072 17208 1106
rect 17242 1072 17258 1106
rect 16643 1020 16650 1060
rect 16333 900 16340 960
rect 16437 927 16487 1007
rect 16643 967 16685 1020
rect 17050 1004 17084 1066
rect 17366 1004 17400 1066
rect 17050 970 17146 1004
rect 17304 970 17400 1004
rect 16634 951 16685 967
rect 16333 871 16349 900
rect 16383 871 16399 900
rect 16437 893 16453 927
rect 16437 877 16487 893
rect 16550 921 16584 944
rect 16333 863 16399 871
rect 16550 825 16584 887
rect 16668 917 16685 951
rect 16634 861 16685 917
rect 14598 791 14627 825
rect 14661 791 14719 825
rect 14753 791 14811 825
rect 14845 791 14903 825
rect 14937 791 14995 825
rect 15029 791 15087 825
rect 15121 791 15179 825
rect 15213 791 15271 825
rect 15305 791 15363 825
rect 15397 791 15455 825
rect 15489 791 15547 825
rect 15581 791 15639 825
rect 15673 791 15731 825
rect 15765 791 15823 825
rect 15857 791 15915 825
rect 15949 791 16007 825
rect 16041 791 16099 825
rect 16133 791 16191 825
rect 16225 791 16283 825
rect 16317 791 16375 825
rect 16409 791 16467 825
rect 16501 791 16559 825
rect 16593 791 16651 825
rect 16685 791 16714 825
rect 17050 814 17146 848
rect 17304 814 17400 848
rect 17050 752 17084 814
rect 17366 752 17400 814
rect 17192 712 17208 746
rect 17242 712 17258 746
rect 17164 662 17198 678
rect 17164 470 17198 486
rect 17252 662 17286 678
rect 17252 470 17286 486
rect 17192 402 17208 436
rect 17242 402 17258 436
rect 17050 334 17084 396
rect 17366 334 17400 396
rect 17050 300 17146 334
rect 17304 300 17400 334
rect 3322 230 3356 292
rect 36 196 132 230
rect 3260 196 3356 230
<< viali >>
rect 8288 5499 9328 5502
rect 8288 5465 9328 5499
rect 8288 5462 9328 5465
rect 840 5257 1000 5260
rect 1960 5257 2120 5260
rect 2740 5257 2900 5260
rect 3660 5257 3820 5260
rect 840 5223 1000 5257
rect 1960 5223 2120 5257
rect 2740 5223 2900 5257
rect 3660 5223 3820 5257
rect 840 5220 1000 5223
rect 1960 5220 2120 5223
rect 2740 5220 2900 5223
rect 3660 5220 3820 5223
rect 1830 5027 1998 5061
rect 2210 5027 2378 5061
rect 2590 5027 3558 5061
rect 3770 5027 3938 5061
rect 1768 4763 1802 4951
rect 2026 4763 2060 4951
rect 2148 4592 2182 4968
rect 2406 4592 2440 4968
rect 2528 4592 2562 4968
rect 3586 4592 3620 4968
rect 3708 4763 3742 4951
rect 3966 4763 4000 4951
rect 1830 4499 1998 4533
rect 2210 4499 2378 4533
rect 2590 4499 3558 4533
rect 3770 4499 3938 4533
rect 450 4347 618 4381
rect 830 4347 998 4381
rect 1088 4347 1256 4381
rect 1470 4347 1638 4381
rect 1728 4347 1896 4381
rect 1986 4347 2154 4381
rect 2244 4347 2412 4381
rect 2630 4347 2798 4381
rect 2888 4347 3056 4381
rect 3146 4347 3314 4381
rect 3404 4347 3572 4381
rect 3790 4347 3958 4381
rect 388 4083 422 4271
rect 646 4083 680 4271
rect 768 3929 802 4117
rect 1026 4083 1060 4271
rect 1284 3929 1318 4117
rect 1408 3929 1442 4117
rect 1666 4083 1700 4271
rect 1924 3929 1958 4117
rect 2182 4083 2216 4271
rect 2440 3929 2474 4117
rect 2568 3929 2602 4117
rect 2826 4083 2860 4271
rect 3084 3929 3118 4117
rect 3342 4083 3376 4271
rect 3600 3929 3634 4117
rect 3728 3929 3762 4117
rect 3986 3929 4020 4117
rect 450 3819 618 3853
rect 830 3819 998 3853
rect 1088 3819 1256 3853
rect 1470 3819 1638 3853
rect 1728 3819 1896 3853
rect 1986 3819 2154 3853
rect 2244 3819 2412 3853
rect 2630 3819 2798 3853
rect 2888 3819 3056 3853
rect 3146 3819 3314 3853
rect 3404 3819 3572 3853
rect 3790 3819 3958 3853
rect 430 3107 598 3141
rect 810 3107 978 3141
rect 1068 3107 1236 3141
rect 1326 3107 1494 3141
rect 1584 3107 1752 3141
rect 1842 3107 2010 3141
rect 2100 3107 2268 3141
rect 2358 3107 2526 3141
rect 2616 3107 2784 3141
rect 2990 3107 3158 3141
rect 368 2843 402 3031
rect 626 2843 660 3031
rect 748 2689 782 2877
rect 1006 2843 1040 3031
rect 1264 2689 1298 2877
rect 1522 2843 1556 3031
rect 1780 2689 1814 2877
rect 2038 2843 2072 3031
rect 2296 2689 2330 2877
rect 2554 2843 2588 3031
rect 2812 2689 2846 2877
rect 2928 2843 2962 3031
rect 3186 2843 3220 3031
rect 3280 2940 3323 3040
rect 3323 2940 3357 3040
rect 3357 2940 3360 3040
rect 430 2579 598 2613
rect 810 2579 978 2613
rect 1068 2579 1236 2613
rect 1326 2579 1494 2613
rect 1584 2579 1752 2613
rect 1842 2579 2010 2613
rect 2100 2579 2268 2613
rect 2358 2579 2526 2613
rect 2616 2579 2784 2613
rect 2990 2579 3158 2613
rect 6096 5329 6264 5363
rect 6354 5329 6522 5363
rect 7256 5329 7424 5363
rect 10208 5329 10376 5363
rect 11096 5329 11264 5363
rect 11354 5329 11522 5363
rect 5776 3765 5810 5253
rect 6034 2311 6068 3799
rect 6292 3765 6326 5253
rect 6550 2311 6584 3799
rect 6808 3765 6842 5253
rect 6936 5111 6970 5199
rect 7194 5165 7228 5253
rect 7452 5111 7486 5199
rect 7710 5165 7744 5253
rect 7968 5111 8002 5199
rect 8226 5165 8260 5253
rect 8484 5111 8518 5199
rect 8742 5165 8776 5253
rect 8856 5111 8890 5199
rect 9114 5165 9148 5253
rect 9372 5111 9406 5199
rect 9630 5165 9664 5253
rect 9888 5111 9922 5199
rect 10146 5165 10180 5253
rect 10404 5111 10438 5199
rect 10662 5165 10696 5253
rect 6998 5001 7166 5035
rect 7256 5001 7424 5035
rect 7514 5001 7682 5035
rect 7772 5001 7940 5035
rect 8030 5001 8198 5035
rect 8288 5001 8456 5035
rect 8546 5001 8714 5035
rect 8938 5001 9086 5035
rect 9086 5001 9106 5035
rect 9196 5001 9344 5035
rect 9344 5001 9364 5035
rect 9454 5001 9602 5035
rect 9602 5001 9622 5035
rect 9712 5001 9860 5035
rect 9860 5001 9880 5035
rect 9970 5001 10118 5035
rect 10118 5001 10138 5035
rect 10208 5001 10376 5035
rect 10466 5001 10634 5035
rect 10634 5001 10654 5035
rect 5838 2201 6006 2235
rect 6612 2201 6780 2235
rect 8784 4648 8818 4682
rect 8976 4648 9010 4682
rect 8640 4339 8674 4477
rect 8736 4443 8770 4581
rect 8832 4339 8866 4477
rect 8928 4443 8962 4581
rect 9024 4339 9058 4477
rect 8688 4238 8722 4272
rect 8880 4238 8914 4272
rect 7682 3928 7850 3962
rect 7940 3928 8108 3962
rect 8198 3928 8366 3962
rect 8456 3928 8624 3962
rect 7620 3719 7654 3807
rect 7878 3773 7912 3861
rect 8136 3719 8170 3807
rect 8394 3773 8428 3861
rect 8842 3868 9010 3902
rect 9100 3868 9268 3902
rect 9358 3868 9526 3902
rect 9616 3868 9784 3902
rect 9874 3868 10042 3902
rect 10132 3868 10300 3902
rect 8652 3719 8686 3807
rect 7682 3618 7850 3652
rect 7940 3618 8108 3652
rect 8198 3618 8366 3652
rect 8456 3618 8624 3652
rect 8780 3313 8814 3801
rect 9038 2859 9072 3347
rect 9296 3313 9330 3801
rect 9554 2859 9588 3347
rect 9812 3313 9846 3801
rect 10070 2859 10104 3347
rect 10328 3313 10362 3801
rect 8842 2758 9010 2792
rect 9100 2758 9268 2792
rect 9358 2758 9526 2792
rect 9616 2758 9784 2792
rect 9874 2758 10042 2792
rect 10132 2758 10300 2792
rect 8108 2652 8208 2682
rect 9528 2652 9628 2682
rect 8108 2618 8208 2652
rect 9528 2618 9628 2652
rect 8108 2602 8208 2618
rect 9528 2602 9628 2618
rect 10776 3765 10810 5253
rect 11034 2311 11068 3799
rect 11292 3765 11326 5253
rect 11550 2311 11584 3799
rect 11808 3765 11842 5253
rect 10838 2201 11006 2235
rect 11612 2201 11780 2235
rect 14566 5337 14604 5734
rect 14732 5337 14770 5734
rect 14898 5337 14936 5734
rect 15064 5337 15102 5734
rect 15230 5337 15268 5734
rect 15396 5337 15434 5734
rect 15562 5337 15600 5734
rect 15728 5337 15766 5734
rect 16040 5337 16078 5734
rect 16206 5337 16244 5734
rect 16372 5337 16410 5734
rect 16538 5337 16576 5734
rect 16704 5337 16742 5734
rect 16870 5337 16908 5734
rect 17036 5337 17074 5734
rect 17202 5337 17240 5734
rect 14566 4006 14604 4403
rect 14732 4006 14770 4403
rect 14898 4006 14936 4403
rect 15064 4006 15102 4403
rect 15230 4006 15268 4403
rect 15396 4006 15434 4403
rect 15562 4006 15600 4403
rect 15728 4006 15766 4403
rect 16040 4006 16078 4403
rect 16206 4006 16244 4403
rect 16372 4006 16410 4403
rect 16538 4006 16576 4403
rect 16704 4006 16742 4403
rect 16870 4006 16908 4403
rect 17036 4006 17074 4403
rect 17202 4006 17240 4403
rect 14616 3169 14654 3566
rect 14782 3169 14820 3566
rect 14948 3169 14986 3566
rect 15114 3169 15152 3566
rect 15280 3169 15318 3566
rect 15446 3169 15484 3566
rect 15612 3169 15650 3566
rect 15778 3169 15816 3566
rect 14616 2338 14654 2735
rect 14782 2338 14820 2735
rect 14948 2338 14986 2735
rect 15114 2338 15152 2735
rect 15280 2338 15318 2735
rect 15446 2338 15484 2735
rect 15612 2338 15650 2735
rect 15778 2338 15816 2735
rect 234 1910 402 1944
rect 614 1910 782 1944
rect 994 1910 1162 1944
rect 1374 1910 1542 1944
rect 1754 1910 1922 1944
rect 2134 1910 2302 1944
rect 2514 1910 2682 1944
rect 2894 1910 3062 1944
rect 172 1684 206 1860
rect 430 1684 464 1860
rect 552 1684 586 1860
rect 810 1684 844 1860
rect 932 1684 966 1860
rect 1190 1684 1224 1860
rect 1312 1684 1346 1860
rect 1570 1684 1604 1860
rect 1692 1684 1726 1860
rect 1950 1684 1984 1860
rect 2072 1684 2106 1860
rect 2330 1684 2364 1860
rect 2452 1684 2486 1860
rect 2710 1684 2744 1860
rect 2832 1684 2866 1860
rect 3090 1684 3124 1860
rect 234 1600 402 1634
rect 614 1600 782 1634
rect 994 1600 1162 1634
rect 1374 1600 1542 1634
rect 1754 1600 1922 1634
rect 2134 1600 2302 1634
rect 2514 1600 2682 1634
rect 2894 1600 3062 1634
rect 234 1492 402 1526
rect 614 1492 782 1526
rect 994 1492 1162 1526
rect 1374 1492 1542 1526
rect 1754 1492 1922 1526
rect 2134 1492 2302 1526
rect 2514 1492 2682 1526
rect 2894 1492 3062 1526
rect 172 1266 206 1442
rect 430 1266 464 1442
rect 552 1266 586 1442
rect 810 1266 844 1442
rect 932 1266 966 1442
rect 1190 1266 1224 1442
rect 1312 1266 1346 1442
rect 1570 1266 1604 1442
rect 1692 1266 1726 1442
rect 1950 1266 1984 1442
rect 2072 1266 2106 1442
rect 2330 1266 2364 1442
rect 2452 1266 2486 1442
rect 2710 1266 2744 1442
rect 2832 1266 2866 1442
rect 3090 1266 3124 1442
rect 234 1182 402 1216
rect 614 1182 782 1216
rect 994 1182 1162 1216
rect 1374 1182 1542 1216
rect 1754 1182 1922 1216
rect 2134 1182 2302 1216
rect 2514 1182 2682 1216
rect 2894 1182 3062 1216
rect 234 1074 402 1108
rect 614 1074 782 1108
rect 994 1074 1162 1108
rect 1374 1074 1542 1108
rect 1754 1074 1922 1108
rect 2134 1074 2302 1108
rect 2514 1074 2682 1108
rect 2894 1074 3062 1108
rect 172 848 206 1024
rect 430 848 464 1024
rect 552 848 586 1024
rect 810 848 844 1024
rect 932 848 966 1024
rect 1190 848 1224 1024
rect 1312 848 1346 1024
rect 1570 848 1604 1024
rect 1692 848 1726 1024
rect 1950 848 1984 1024
rect 2072 848 2106 1024
rect 2330 848 2364 1024
rect 2452 848 2486 1024
rect 2710 848 2744 1024
rect 2832 848 2866 1024
rect 3090 848 3124 1024
rect 234 764 402 798
rect 614 764 782 798
rect 994 764 1162 798
rect 1374 764 1542 798
rect 1754 764 1922 798
rect 2134 764 2302 798
rect 2514 764 2682 798
rect 2894 764 3062 798
rect 234 656 402 690
rect 614 656 782 690
rect 994 656 1162 690
rect 1374 656 1542 690
rect 1754 656 1922 690
rect 2134 656 2302 690
rect 2514 656 2682 690
rect 2894 656 3062 690
rect 172 430 206 606
rect 430 430 464 606
rect 552 430 586 606
rect 810 430 844 606
rect 932 430 966 606
rect 1190 430 1224 606
rect 1312 430 1346 606
rect 1570 430 1604 606
rect 1692 430 1726 606
rect 1950 430 1984 606
rect 2072 430 2106 606
rect 2330 430 2364 606
rect 2452 430 2486 606
rect 2710 430 2744 606
rect 2832 430 2866 606
rect 3090 430 3124 606
rect 234 346 402 380
rect 614 346 782 380
rect 994 346 1162 380
rect 1374 346 1542 380
rect 1754 346 1922 380
rect 2134 346 2302 380
rect 2514 346 2682 380
rect 2894 346 3062 380
rect 14627 1335 14661 1369
rect 14719 1335 14753 1369
rect 14811 1335 14845 1369
rect 14903 1335 14937 1369
rect 14995 1335 15029 1369
rect 15087 1335 15121 1369
rect 15179 1335 15213 1369
rect 15271 1335 15305 1369
rect 15363 1335 15397 1369
rect 15455 1335 15489 1369
rect 15547 1335 15581 1369
rect 15639 1335 15673 1369
rect 15731 1335 15765 1369
rect 15823 1335 15857 1369
rect 15915 1335 15949 1369
rect 16007 1335 16041 1369
rect 16099 1335 16133 1369
rect 16191 1335 16225 1369
rect 16283 1335 16317 1369
rect 16375 1335 16409 1369
rect 16467 1335 16501 1369
rect 16559 1335 16593 1369
rect 16651 1335 16685 1369
rect 14430 1290 14500 1300
rect 14430 1250 14450 1290
rect 14450 1250 14490 1290
rect 14490 1250 14500 1290
rect 14620 1057 14660 1080
rect 14620 1023 14630 1057
rect 14630 1023 14660 1057
rect 14620 1020 14660 1023
rect 14720 1038 14732 1063
rect 14732 1038 14754 1063
rect 14720 1029 14754 1038
rect 14801 1183 14835 1199
rect 14801 1165 14835 1183
rect 14900 950 14960 990
rect 15179 1165 15213 1199
rect 15087 1029 15121 1063
rect 15803 1173 15837 1199
rect 15803 1165 15834 1173
rect 15834 1165 15837 1173
rect 15359 961 15393 995
rect 15431 977 15455 995
rect 15455 977 15465 995
rect 15431 961 15465 977
rect 15803 1047 15837 1063
rect 15803 1029 15829 1047
rect 15829 1029 15837 1047
rect 16019 1049 16053 1058
rect 16019 1024 16035 1049
rect 16035 1024 16053 1049
rect 16079 961 16113 995
rect 17208 1800 17242 1834
rect 17164 1165 17198 1741
rect 17252 1165 17286 1741
rect 17360 1180 17366 1740
rect 17366 1180 17400 1740
rect 17208 1072 17242 1106
rect 16650 1020 16690 1060
rect 16340 939 16349 960
rect 16349 939 16383 960
rect 16383 939 16400 960
rect 16340 905 16400 939
rect 16340 900 16349 905
rect 16349 900 16383 905
rect 16383 900 16400 905
rect 14627 791 14661 825
rect 14719 791 14753 825
rect 14811 791 14845 825
rect 14903 791 14937 825
rect 14995 791 15029 825
rect 15087 791 15121 825
rect 15179 791 15213 825
rect 15271 791 15305 825
rect 15363 791 15397 825
rect 15455 791 15489 825
rect 15547 791 15581 825
rect 15639 791 15673 825
rect 15731 791 15765 825
rect 15823 791 15857 825
rect 15915 791 15949 825
rect 16007 791 16041 825
rect 16099 791 16133 825
rect 16191 791 16225 825
rect 16283 791 16317 825
rect 16375 791 16409 825
rect 16467 791 16501 825
rect 16559 791 16593 825
rect 16651 791 16685 825
rect 17208 712 17242 746
rect 17164 486 17198 662
rect 17252 486 17286 662
rect 17360 480 17366 640
rect 17366 480 17400 640
rect 17208 402 17242 436
rect 220 230 440 240
rect 1100 230 1320 240
rect 2020 230 2240 240
rect 2860 230 3080 240
rect 220 200 440 230
rect 1100 200 1320 230
rect 2020 200 2240 230
rect 2860 200 3080 230
<< metal1 >>
rect 6940 7200 7260 7540
rect 6900 7160 7300 7200
rect 6900 6880 6940 7160
rect 7260 6880 7300 7160
rect 6900 6860 7300 6880
rect 200 6760 13100 6780
rect 200 6580 12880 6760
rect 590 6560 12880 6580
rect 13080 6560 13100 6760
rect 8750 5742 8760 5900
rect 320 5480 4240 5500
rect 320 5400 3500 5480
rect 310 5300 320 5400
rect 400 5300 1600 5400
rect 1720 5320 3500 5400
rect 4000 5400 4240 5480
rect 6268 5442 6288 5562
rect 6348 5542 8468 5562
rect 8748 5542 8760 5742
rect 6348 5442 8188 5542
rect 8288 5540 8760 5542
rect 8960 5542 8970 5900
rect 14560 5740 14610 5746
rect 14726 5740 14776 5746
rect 14540 5734 14776 5740
rect 8960 5540 9328 5542
rect 8288 5502 9328 5540
rect 8288 5442 9328 5462
rect 9428 5522 11368 5542
rect 9428 5442 11268 5522
rect 6268 5422 11268 5442
rect 11328 5422 11368 5522
rect 4000 5320 4040 5400
rect 1720 5300 4040 5320
rect 4140 5300 4240 5400
rect 12020 5400 14480 5420
rect 6084 5363 6276 5369
rect 6084 5362 6096 5363
rect 5828 5329 6096 5362
rect 6264 5362 6276 5363
rect 6342 5363 6534 5369
rect 6342 5362 6354 5363
rect 6264 5329 6354 5362
rect 6522 5362 6534 5363
rect 7244 5363 7436 5369
rect 7244 5362 7256 5363
rect 6522 5329 7256 5362
rect 7424 5329 7436 5363
rect 5828 5323 7436 5329
rect 10188 5363 11788 5382
rect 10188 5329 10208 5363
rect 10376 5329 11096 5363
rect 11264 5329 11354 5363
rect 11522 5329 11788 5363
rect 5828 5322 7428 5323
rect 10188 5322 11788 5329
rect 840 5266 1000 5300
rect 1960 5266 2120 5300
rect 2740 5266 2900 5300
rect 3660 5266 3820 5300
rect 828 5260 1012 5266
rect 828 5220 840 5260
rect 1000 5220 1012 5260
rect 828 5214 1012 5220
rect 1948 5260 2132 5266
rect 1948 5220 1960 5260
rect 2120 5220 2132 5260
rect 1948 5214 2132 5220
rect 2728 5260 2912 5266
rect 2728 5220 2740 5260
rect 2900 5220 2912 5260
rect 2728 5214 2912 5220
rect 3648 5260 3832 5266
rect 3648 5220 3660 5260
rect 3820 5220 3832 5260
rect 3648 5214 3832 5220
rect 5770 5253 5816 5265
rect 1820 5067 2040 5080
rect 1818 5061 2040 5067
rect 1818 5060 1830 5061
rect 1800 5027 1830 5060
rect 1998 5027 2040 5061
rect 1800 4963 2040 5027
rect 2198 5061 2390 5067
rect 2198 5027 2210 5061
rect 2378 5027 2390 5061
rect 2198 5021 2390 5027
rect 2578 5061 3570 5067
rect 2578 5027 2590 5061
rect 3558 5027 3570 5061
rect 3758 5061 3950 5067
rect 3758 5040 3770 5061
rect 2578 5021 3570 5027
rect 3720 5027 3770 5040
rect 3938 5060 3950 5061
rect 3938 5027 3980 5060
rect 2142 4968 2188 4980
rect 1762 4960 2066 4963
rect 2142 4960 2148 4968
rect 1590 4840 1600 4960
rect 1720 4951 2148 4960
rect 1720 4840 1768 4951
rect 1762 4763 1768 4840
rect 1802 4840 2026 4951
rect 1802 4763 1808 4840
rect 1762 4751 1808 4763
rect 2020 4763 2026 4840
rect 2060 4840 2148 4951
rect 2060 4763 2066 4840
rect 2020 4751 2066 4763
rect 2142 4592 2148 4840
rect 2182 4960 2188 4968
rect 2400 4968 2446 4980
rect 2182 4840 2200 4960
rect 2182 4592 2188 4840
rect 2400 4800 2406 4968
rect 2440 4800 2446 4968
rect 2522 4968 2568 4980
rect 2142 4580 2188 4592
rect 2350 4580 2360 4800
rect 2440 4580 2450 4800
rect 2522 4760 2528 4968
rect 2520 4620 2528 4760
rect 2522 4592 2528 4620
rect 2562 4760 2568 4968
rect 3580 4968 3626 4980
rect 2562 4740 3380 4760
rect 2562 4620 3280 4740
rect 3380 4620 3390 4740
rect 2562 4592 2568 4620
rect 2522 4580 2568 4592
rect 3580 4592 3586 4968
rect 3620 4960 3626 4968
rect 3720 4963 3980 5027
rect 3702 4960 4006 4963
rect 3620 4951 4040 4960
rect 3620 4820 3708 4951
rect 3620 4592 3626 4820
rect 3702 4763 3708 4820
rect 3742 4820 3966 4951
rect 3742 4763 3748 4820
rect 3702 4751 3748 4763
rect 3960 4763 3966 4820
rect 4000 4840 4040 4951
rect 4140 4840 4150 4960
rect 4000 4820 4020 4840
rect 4000 4763 4006 4820
rect 3960 4751 4006 4763
rect 3580 4580 3626 4592
rect 2200 4539 2620 4540
rect 1818 4533 2010 4539
rect 1818 4499 1830 4533
rect 1998 4499 2010 4533
rect 1818 4493 2010 4499
rect 2198 4533 2620 4539
rect 2720 4539 2730 4540
rect 2720 4533 3570 4539
rect 2198 4499 2210 4533
rect 2378 4500 2590 4533
rect 2378 4499 2390 4500
rect 2198 4493 2390 4499
rect 2578 4499 2590 4500
rect 3558 4499 3570 4533
rect 2578 4493 2620 4499
rect 2610 4480 2620 4493
rect 2720 4493 3570 4499
rect 3758 4533 3950 4539
rect 3758 4499 3770 4533
rect 3938 4499 3950 4533
rect 3758 4493 3950 4499
rect 2720 4480 2730 4493
rect 438 4381 630 4387
rect 438 4347 450 4381
rect 618 4380 630 4381
rect 818 4381 1010 4387
rect 618 4347 640 4380
rect 438 4341 640 4347
rect 818 4347 830 4381
rect 998 4347 1010 4381
rect 818 4341 1010 4347
rect 1076 4381 1268 4387
rect 1076 4347 1088 4381
rect 1256 4347 1268 4381
rect 1076 4341 1268 4347
rect 1458 4381 1650 4387
rect 1458 4347 1470 4381
rect 1638 4347 1650 4381
rect 1458 4341 1650 4347
rect 1716 4381 1908 4387
rect 1716 4347 1728 4381
rect 1896 4347 1908 4381
rect 1716 4341 1908 4347
rect 1974 4381 2166 4387
rect 1974 4347 1986 4381
rect 2154 4347 2166 4381
rect 1974 4341 2166 4347
rect 2232 4381 2424 4387
rect 2232 4347 2244 4381
rect 2412 4347 2424 4381
rect 2232 4341 2424 4347
rect 2618 4381 2810 4387
rect 2618 4347 2630 4381
rect 2798 4347 2810 4381
rect 2618 4341 2810 4347
rect 2876 4381 3068 4387
rect 2876 4347 2888 4381
rect 3056 4347 3068 4381
rect 2876 4341 3068 4347
rect 3134 4381 3326 4387
rect 3134 4347 3146 4381
rect 3314 4347 3326 4381
rect 3134 4341 3326 4347
rect 3392 4381 3584 4387
rect 3392 4347 3404 4381
rect 3572 4347 3584 4381
rect 3392 4341 3584 4347
rect 3778 4381 3970 4387
rect 3778 4347 3790 4381
rect 3958 4347 3970 4381
rect 3778 4341 3970 4347
rect 440 4300 640 4341
rect 310 4220 320 4300
rect 400 4283 1060 4300
rect 400 4271 1066 4283
rect 422 4220 646 4271
rect 382 4083 388 4220
rect 422 4083 428 4220
rect 382 4071 428 4083
rect 640 4083 646 4220
rect 680 4220 1026 4271
rect 680 4083 686 4220
rect 640 4071 686 4083
rect 762 4117 808 4129
rect 762 4020 768 4117
rect 760 3929 768 4020
rect 802 4020 808 4117
rect 1020 4083 1026 4220
rect 1060 4083 1066 4271
rect 1660 4271 2360 4300
rect 1020 4071 1066 4083
rect 1278 4117 1324 4129
rect 1278 4020 1284 4117
rect 802 3929 1284 4020
rect 1318 3929 1324 4117
rect 1402 4117 1448 4129
rect 1402 4000 1408 4117
rect 760 3917 1324 3929
rect 1400 3929 1408 4000
rect 1442 4000 1448 4117
rect 1660 4083 1666 4271
rect 1700 4200 2182 4271
rect 1700 4083 1706 4200
rect 1660 4071 1706 4083
rect 1918 4117 1964 4129
rect 1918 4000 1924 4117
rect 1442 3929 1924 4000
rect 1958 4000 1964 4117
rect 2176 4083 2182 4200
rect 2216 4200 2360 4271
rect 2440 4200 2500 4300
rect 2820 4280 2866 4283
rect 3336 4280 3382 4283
rect 2820 4271 2920 4280
rect 2216 4083 2222 4200
rect 2176 4071 2222 4083
rect 2434 4117 2480 4129
rect 2434 4000 2440 4117
rect 1958 3929 2440 4000
rect 2474 4000 2480 4117
rect 2562 4117 2608 4129
rect 2562 4000 2568 4117
rect 2474 3929 2568 4000
rect 2602 4000 2608 4117
rect 2820 4083 2826 4271
rect 2860 4180 2920 4271
rect 3020 4271 3382 4280
rect 3020 4180 3342 4271
rect 2860 4083 2866 4180
rect 2820 4071 2866 4083
rect 3078 4117 3124 4129
rect 3078 4000 3084 4117
rect 2602 3929 3084 4000
rect 3118 4000 3124 4117
rect 3336 4083 3342 4180
rect 3376 4083 3382 4271
rect 3336 4071 3382 4083
rect 3594 4117 3640 4129
rect 3594 4000 3600 4117
rect 3118 3929 3600 4000
rect 3634 4000 3640 4117
rect 3722 4117 3768 4129
rect 3722 4000 3728 4117
rect 3634 3929 3728 4000
rect 3762 4000 3768 4117
rect 3980 4117 4026 4129
rect 3980 4000 3986 4117
rect 3762 3929 3986 4000
rect 4020 4000 4026 4117
rect 4020 3929 4040 4000
rect 760 3860 1320 3917
rect 1400 3900 4040 3929
rect 438 3853 630 3859
rect 438 3819 450 3853
rect 618 3819 630 3853
rect 760 3853 840 3860
rect 940 3859 2420 3860
rect 940 3853 2424 3859
rect 760 3840 830 3853
rect 438 3813 630 3819
rect 818 3819 830 3840
rect 998 3819 1088 3853
rect 1256 3819 1470 3853
rect 1638 3819 1728 3853
rect 1896 3819 1986 3853
rect 2154 3819 2244 3853
rect 2412 3819 2424 3853
rect 818 3813 840 3819
rect 820 3800 840 3813
rect 940 3813 2424 3819
rect 940 3800 2420 3813
rect 2610 3800 2620 3860
rect 2720 3859 3580 3860
rect 3780 3859 3960 3900
rect 5770 3862 5776 5253
rect 2720 3853 3584 3859
rect 2798 3820 2888 3853
rect 2798 3819 2810 3820
rect 2720 3813 2810 3819
rect 2876 3819 2888 3820
rect 3056 3820 3146 3853
rect 3056 3819 3068 3820
rect 2876 3813 3068 3819
rect 3134 3819 3146 3820
rect 3314 3820 3404 3853
rect 3314 3819 3326 3820
rect 3134 3813 3326 3819
rect 3392 3819 3404 3820
rect 3572 3819 3584 3853
rect 3392 3813 3584 3819
rect 3778 3853 3970 3859
rect 3778 3819 3790 3853
rect 3958 3819 3970 3853
rect 3778 3813 3970 3819
rect 2720 3800 2730 3813
rect 5768 3765 5776 3862
rect 5810 3862 5816 5253
rect 6286 5253 6332 5265
rect 6286 5122 6292 5253
rect 6326 5122 6332 5253
rect 6802 5253 6848 5265
rect 6258 4882 6268 5122
rect 6368 4882 6378 5122
rect 5810 3811 6048 3862
rect 5810 3799 6074 3811
rect 5810 3765 6034 3799
rect 5768 3682 6034 3765
rect 4040 3540 4370 3560
rect 2610 3420 2620 3540
rect 2720 3420 4370 3540
rect 2620 3400 4370 3420
rect 4040 3360 4370 3400
rect 380 3141 640 3160
rect 380 3107 430 3141
rect 598 3107 640 3141
rect 380 3043 640 3107
rect 798 3141 990 3147
rect 798 3107 810 3141
rect 978 3107 990 3141
rect 798 3101 990 3107
rect 1056 3141 1248 3147
rect 1056 3107 1068 3141
rect 1236 3107 1248 3141
rect 1056 3101 1248 3107
rect 1314 3141 1506 3147
rect 1314 3107 1326 3141
rect 1494 3107 1506 3141
rect 1314 3101 1506 3107
rect 1572 3141 1764 3147
rect 1572 3107 1584 3141
rect 1752 3107 1764 3141
rect 1572 3101 1764 3107
rect 1830 3141 2022 3147
rect 1830 3107 1842 3141
rect 2010 3107 2022 3141
rect 1830 3101 2022 3107
rect 2088 3141 2280 3147
rect 2088 3107 2100 3141
rect 2268 3107 2280 3141
rect 2088 3101 2280 3107
rect 2346 3141 2538 3147
rect 2346 3107 2358 3141
rect 2526 3107 2538 3141
rect 2346 3101 2538 3107
rect 2604 3141 2796 3147
rect 2604 3107 2616 3141
rect 2784 3107 2796 3141
rect 2604 3101 2796 3107
rect 2960 3141 3180 3160
rect 2960 3107 2990 3141
rect 3158 3107 3180 3141
rect 2960 3043 3180 3107
rect 362 3040 666 3043
rect 1000 3040 1046 3043
rect 1516 3040 1562 3043
rect 2032 3040 2078 3043
rect 2548 3040 2594 3043
rect 2922 3040 3226 3043
rect 3274 3040 3366 3052
rect 4040 3040 4380 3100
rect 360 3031 3280 3040
rect 360 2940 368 3031
rect 362 2843 368 2940
rect 402 2940 626 3031
rect 402 2843 408 2940
rect 362 2831 408 2843
rect 620 2843 626 2940
rect 660 2940 1006 3031
rect 660 2843 666 2940
rect 620 2831 666 2843
rect 742 2877 788 2889
rect 742 2800 748 2877
rect 740 2689 748 2800
rect 782 2800 788 2877
rect 1000 2843 1006 2940
rect 1040 2940 1522 3031
rect 1040 2843 1046 2940
rect 1000 2831 1046 2843
rect 1258 2877 1304 2889
rect 1258 2800 1264 2877
rect 782 2689 1264 2800
rect 1298 2800 1304 2877
rect 1516 2843 1522 2940
rect 1556 2940 2038 3031
rect 1556 2843 1562 2940
rect 1516 2831 1562 2843
rect 1774 2877 1820 2889
rect 1774 2800 1780 2877
rect 1298 2689 1780 2800
rect 1814 2800 1820 2877
rect 2032 2843 2038 2940
rect 2072 2940 2554 3031
rect 2072 2843 2078 2940
rect 2032 2831 2078 2843
rect 2290 2877 2336 2889
rect 2290 2800 2296 2877
rect 1814 2689 2296 2800
rect 2330 2800 2336 2877
rect 2548 2843 2554 2940
rect 2588 2940 2928 3031
rect 2588 2843 2594 2940
rect 2548 2831 2594 2843
rect 2806 2877 2852 2889
rect 2806 2800 2812 2877
rect 2330 2780 2812 2800
rect 2330 2689 2620 2780
rect 418 2613 610 2619
rect 418 2579 430 2613
rect 598 2579 610 2613
rect 418 2573 610 2579
rect 740 2613 2620 2689
rect 2700 2689 2812 2780
rect 2846 2689 2852 2877
rect 2922 2843 2928 2940
rect 2962 2940 3186 3031
rect 2962 2843 2968 2940
rect 2922 2831 2968 2843
rect 3180 2843 3186 2940
rect 3220 2940 3280 3031
rect 3400 2940 4380 3040
rect 3220 2843 3226 2940
rect 3274 2928 3366 2940
rect 4040 2900 4380 2940
rect 4560 3080 5560 3100
rect 4560 2920 5380 3080
rect 5540 2920 5560 3080
rect 4560 2900 5560 2920
rect 3180 2831 3226 2843
rect 2700 2677 2852 2689
rect 2700 2613 2840 2677
rect 740 2579 810 2613
rect 978 2579 1068 2613
rect 1236 2579 1326 2613
rect 1494 2579 1584 2613
rect 1752 2579 1842 2613
rect 2010 2579 2100 2613
rect 2268 2579 2358 2613
rect 2526 2579 2616 2613
rect 2784 2579 2840 2613
rect 740 2560 2840 2579
rect 2978 2613 3170 2619
rect 2978 2579 2990 2613
rect 3158 2579 3170 2613
rect 2978 2573 3170 2579
rect 2030 2420 2040 2480
rect 2100 2420 2920 2480
rect 3020 2420 3030 2480
rect 530 2240 540 2320
rect 600 2300 1180 2320
rect 600 2240 840 2300
rect 940 2240 1180 2300
rect 1240 2240 1250 2320
rect 1290 2280 1300 2360
rect 1360 2280 1940 2360
rect 2000 2280 2620 2360
rect 2720 2280 2730 2360
rect 6028 2311 6034 3682
rect 6068 3142 6074 3799
rect 6286 3765 6292 4882
rect 6326 3765 6332 4882
rect 6802 3862 6808 5253
rect 6548 3811 6808 3862
rect 6286 3753 6332 3765
rect 6544 3799 6808 3811
rect 6544 3142 6550 3799
rect 6068 3042 6550 3142
rect 6068 2542 6074 3042
rect 6068 2311 6088 2542
rect 6028 2242 6088 2311
rect 6544 2311 6550 3042
rect 6584 3765 6808 3799
rect 6842 3765 6848 5253
rect 7188 5253 8188 5282
rect 7188 5242 7194 5253
rect 6948 5211 7194 5242
rect 6930 5199 7194 5211
rect 6930 5111 6936 5199
rect 6970 5165 7194 5199
rect 7228 5242 7710 5253
rect 7228 5165 7234 5242
rect 6970 5153 7234 5165
rect 7446 5199 7492 5211
rect 6970 5111 7208 5153
rect 7446 5122 7452 5199
rect 6930 5099 7208 5111
rect 6948 5035 7208 5099
rect 7428 5111 7452 5122
rect 7486 5122 7492 5199
rect 7704 5165 7710 5242
rect 7744 5242 8188 5253
rect 7744 5165 7750 5242
rect 7704 5153 7750 5165
rect 7962 5199 8008 5211
rect 8178 5202 8188 5242
rect 8288 5202 8298 5282
rect 8508 5265 8768 5282
rect 9128 5265 10188 5282
rect 8508 5253 8782 5265
rect 8508 5211 8742 5253
rect 7962 5122 7968 5199
rect 7486 5111 7968 5122
rect 8002 5122 8008 5199
rect 8220 5165 8226 5202
rect 8260 5165 8266 5202
rect 8478 5199 8742 5211
rect 8478 5182 8484 5199
rect 8518 5182 8742 5199
rect 8220 5153 8266 5165
rect 8458 5122 8468 5182
rect 8002 5111 8468 5122
rect 8548 5165 8742 5182
rect 8776 5165 8782 5253
rect 9108 5253 10188 5265
rect 10656 5262 10702 5265
rect 9108 5242 9114 5253
rect 9148 5242 9630 5253
rect 8888 5211 9108 5242
rect 8548 5153 8782 5165
rect 8850 5199 9108 5211
rect 7428 5082 8468 5111
rect 8548 5082 8768 5153
rect 8850 5111 8856 5199
rect 8890 5162 9108 5199
rect 9188 5162 9198 5242
rect 9366 5202 9412 5211
rect 8890 5153 9154 5162
rect 8890 5111 9148 5153
rect 8850 5102 9148 5111
rect 8850 5099 9208 5102
rect 8268 5042 8468 5082
rect 7248 5041 8468 5042
rect 6948 5002 6998 5035
rect 6986 5001 6998 5002
rect 7166 5002 7208 5035
rect 7244 5035 8468 5041
rect 7166 5001 7178 5002
rect 6986 4995 7178 5001
rect 7244 5001 7256 5035
rect 7424 5002 7514 5035
rect 7424 5001 7436 5002
rect 7244 4995 7436 5001
rect 7502 5001 7514 5002
rect 7682 5002 7772 5035
rect 7682 5001 7694 5002
rect 7502 4995 7694 5001
rect 7760 5001 7772 5002
rect 7940 5002 8030 5035
rect 7940 5001 7952 5002
rect 7760 4995 7952 5001
rect 8018 5001 8030 5002
rect 8198 5002 8288 5035
rect 8198 5001 8210 5002
rect 8018 4995 8210 5001
rect 8276 5001 8288 5002
rect 8456 5001 8468 5035
rect 8508 5035 8768 5082
rect 8508 5002 8546 5035
rect 8276 4995 8468 5001
rect 8534 5001 8546 5002
rect 8714 5002 8768 5035
rect 8888 5042 9208 5099
rect 9338 5082 9348 5202
rect 9428 5122 9438 5202
rect 9624 5165 9630 5242
rect 9664 5242 10146 5253
rect 9664 5165 9670 5242
rect 9624 5153 9670 5165
rect 9882 5199 9928 5211
rect 9882 5122 9888 5199
rect 9428 5111 9888 5122
rect 9922 5122 9928 5199
rect 10140 5165 10146 5242
rect 10180 5242 10188 5253
rect 10548 5253 10708 5262
rect 10180 5165 10186 5242
rect 10140 5153 10186 5165
rect 10398 5202 10444 5211
rect 10548 5202 10662 5253
rect 10398 5199 10662 5202
rect 10398 5122 10404 5199
rect 9922 5111 10404 5122
rect 10438 5165 10662 5199
rect 10696 5165 10708 5253
rect 10438 5162 10708 5165
rect 10770 5253 10816 5265
rect 10438 5153 10702 5162
rect 10438 5111 10688 5153
rect 9428 5082 10688 5111
rect 8888 5041 10368 5042
rect 8888 5035 10388 5041
rect 8888 5002 8938 5035
rect 8714 5001 8726 5002
rect 8534 4995 8726 5001
rect 8926 5001 8938 5002
rect 9106 5002 9196 5035
rect 9106 5001 9118 5002
rect 8926 4995 9118 5001
rect 9184 5001 9196 5002
rect 9364 5002 9454 5035
rect 9364 5001 9376 5002
rect 9184 4995 9376 5001
rect 9442 5001 9454 5002
rect 9622 5002 9712 5035
rect 9622 5001 9634 5002
rect 9442 4995 9634 5001
rect 9700 5001 9712 5002
rect 9880 5002 9970 5035
rect 9880 5001 9892 5002
rect 9700 4995 9892 5001
rect 9958 5001 9970 5002
rect 10138 5002 10208 5035
rect 10138 5001 10150 5002
rect 9958 4995 10150 5001
rect 10196 5001 10208 5002
rect 10376 5001 10388 5035
rect 10448 5035 10688 5082
rect 10448 5022 10466 5035
rect 10196 4995 10388 5001
rect 10454 5001 10466 5022
rect 10654 5002 10688 5035
rect 10654 5001 10666 5002
rect 10454 4995 10666 5001
rect 8758 4742 8768 4822
rect 8848 4742 10528 4822
rect 10608 4742 10618 4822
rect 8758 4642 8768 4702
rect 8848 4642 8858 4702
rect 8968 4688 9028 4702
rect 8964 4682 9028 4688
rect 8964 4662 8976 4682
rect 8948 4648 8976 4662
rect 9010 4662 9028 4682
rect 9010 4648 9048 4662
rect 8948 4602 9048 4648
rect 8458 4522 8468 4602
rect 8548 4593 8748 4602
rect 8948 4593 9108 4602
rect 8548 4581 8776 4593
rect 8548 4522 8736 4581
rect 8628 4477 8736 4522
rect 8628 4339 8640 4477
rect 8674 4443 8736 4477
rect 8770 4443 8776 4581
rect 8922 4581 9108 4593
rect 8674 4431 8776 4443
rect 8826 4477 8872 4489
rect 8674 4339 8748 4431
rect 8826 4402 8832 4477
rect 8866 4402 8872 4477
rect 8922 4443 8928 4581
rect 8962 4522 9108 4581
rect 9188 4522 9198 4602
rect 8962 4489 9048 4522
rect 8962 4477 9064 4489
rect 8962 4443 9024 4477
rect 8922 4431 9024 4443
rect 8628 4322 8748 4339
rect 8798 4322 8808 4402
rect 8868 4322 8878 4402
rect 8948 4382 9024 4431
rect 9018 4339 9024 4382
rect 9058 4339 9064 4477
rect 9018 4327 9064 4339
rect 8668 4272 8748 4322
rect 8668 4238 8688 4272
rect 8722 4238 8748 4272
rect 8668 4222 8748 4238
rect 8868 4272 8928 4282
rect 8868 4238 8880 4272
rect 8914 4262 8928 4272
rect 9098 4262 9108 4282
rect 8914 4238 9108 4262
rect 8868 4222 9108 4238
rect 9168 4262 9178 4282
rect 9168 4222 9188 4262
rect 7038 4102 7048 4162
rect 7108 4102 9108 4162
rect 9168 4102 9188 4162
rect 8378 4002 8388 4062
rect 8468 4002 8808 4062
rect 8868 4002 8878 4062
rect 7670 3962 7862 3968
rect 7670 3928 7682 3962
rect 7850 3928 7862 3962
rect 7670 3922 7862 3928
rect 7928 3962 8120 3968
rect 7928 3928 7940 3962
rect 8108 3928 8120 3962
rect 7928 3922 8120 3928
rect 8186 3962 8378 3968
rect 8186 3928 8198 3962
rect 8366 3928 8378 3962
rect 8186 3922 8378 3928
rect 8444 3962 8636 3968
rect 8444 3928 8456 3962
rect 8624 3928 8668 3962
rect 8444 3922 8668 3928
rect 7688 3822 7828 3922
rect 8468 3882 8668 3922
rect 9108 3908 10048 3922
rect 8830 3902 9022 3908
rect 8408 3873 8668 3882
rect 7872 3861 7918 3873
rect 8388 3862 8668 3873
rect 7872 3822 7878 3861
rect 7912 3822 7918 3861
rect 6584 3753 6848 3765
rect 7608 3807 7878 3822
rect 6584 3682 6828 3753
rect 7608 3742 7620 3807
rect 7614 3719 7620 3742
rect 7654 3773 7878 3807
rect 7654 3742 7908 3773
rect 7988 3742 7998 3822
rect 8130 3807 8176 3819
rect 8130 3802 8136 3807
rect 8170 3802 8176 3807
rect 7654 3719 7660 3742
rect 7614 3707 7660 3719
rect 6584 3142 6590 3682
rect 7688 3658 7828 3742
rect 7908 3662 7988 3742
rect 8098 3702 8108 3802
rect 8208 3702 8218 3802
rect 8378 3762 8388 3862
rect 8448 3819 8668 3862
rect 8788 3868 8842 3902
rect 9010 3868 9022 3902
rect 8788 3862 9022 3868
rect 9088 3902 10054 3908
rect 9088 3868 9100 3902
rect 9268 3868 9358 3902
rect 9526 3868 9616 3902
rect 9784 3868 9874 3902
rect 10042 3868 10054 3902
rect 9088 3862 10054 3868
rect 10120 3902 10312 3908
rect 10120 3868 10132 3902
rect 10300 3868 10348 3902
rect 10120 3862 10348 3868
rect 8448 3807 8692 3819
rect 8788 3813 9008 3862
rect 8448 3762 8652 3807
rect 8388 3761 8652 3762
rect 8408 3742 8652 3761
rect 8468 3719 8652 3742
rect 8686 3719 8692 3807
rect 8468 3707 8692 3719
rect 8774 3801 9008 3813
rect 7670 3652 7862 3658
rect 7670 3618 7682 3652
rect 7850 3618 7862 3652
rect 7908 3652 8388 3662
rect 8468 3658 8668 3707
rect 7908 3622 7940 3652
rect 7670 3612 7862 3618
rect 7928 3618 7940 3622
rect 8108 3622 8198 3652
rect 8108 3618 8120 3622
rect 7928 3612 8120 3618
rect 8186 3618 8198 3622
rect 8366 3622 8388 3652
rect 8444 3652 8668 3658
rect 8366 3618 8378 3622
rect 8186 3612 8378 3618
rect 8444 3618 8456 3652
rect 8624 3622 8668 3652
rect 8624 3618 8636 3622
rect 8444 3612 8636 3618
rect 8774 3362 8780 3801
rect 8768 3313 8780 3362
rect 8814 3762 9008 3801
rect 9108 3813 9308 3862
rect 10128 3813 10348 3862
rect 10770 3842 10776 5253
rect 9108 3802 9336 3813
rect 8814 3362 8820 3762
rect 9108 3702 9148 3802
rect 8848 3682 9148 3702
rect 8848 3622 8868 3682
rect 8928 3622 9148 3682
rect 9208 3801 9336 3802
rect 9208 3622 9296 3801
rect 8848 3602 9296 3622
rect 8814 3359 9068 3362
rect 8814 3347 9078 3359
rect 8814 3313 9038 3347
rect 8768 3242 9038 3313
rect 6584 3122 8938 3142
rect 6584 3062 8868 3122
rect 8928 3062 8938 3122
rect 6584 3042 8938 3062
rect 6584 2542 6590 3042
rect 9032 2942 9038 3242
rect 8828 2859 9038 2942
rect 9072 3122 9078 3347
rect 9290 3313 9296 3602
rect 9330 3313 9336 3801
rect 9806 3801 9852 3813
rect 9290 3301 9336 3313
rect 9548 3347 9594 3359
rect 9548 3122 9554 3347
rect 9072 3102 9554 3122
rect 9588 3122 9594 3347
rect 9806 3313 9812 3801
rect 9846 3582 9852 3801
rect 10128 3801 10368 3813
rect 10128 3722 10328 3801
rect 9846 3562 10268 3582
rect 9846 3502 10188 3562
rect 10248 3502 10268 3562
rect 9846 3482 10268 3502
rect 9846 3313 9852 3482
rect 10322 3362 10328 3722
rect 10068 3359 10328 3362
rect 9806 3301 9852 3313
rect 10064 3347 10328 3359
rect 10064 3122 10070 3347
rect 9072 3022 9528 3102
rect 9072 2859 9078 3022
rect 9518 2862 9528 3022
rect 9588 3022 10070 3122
rect 9588 2862 9598 3022
rect 8828 2847 9078 2859
rect 9548 2859 9554 2862
rect 9588 2859 9594 2862
rect 9548 2847 9594 2859
rect 10064 2859 10070 3022
rect 10104 3313 10328 3347
rect 10362 3313 10368 3801
rect 10768 3765 10776 3842
rect 10810 3842 10816 5253
rect 11286 5253 11332 5265
rect 11286 5242 11292 5253
rect 11326 5242 11332 5253
rect 11802 5253 11848 5265
rect 11258 4682 11268 5242
rect 11328 4682 11338 5242
rect 10810 3811 11068 3842
rect 10810 3799 11074 3811
rect 10810 3765 11034 3799
rect 10768 3662 11034 3765
rect 10104 3302 10368 3313
rect 10104 2902 10110 3302
rect 10322 3301 10368 3302
rect 11028 3202 11034 3662
rect 10208 3182 10528 3202
rect 10198 3122 10208 3182
rect 10268 3142 10528 3182
rect 10588 3142 11034 3202
rect 10268 3122 11034 3142
rect 10104 2859 10268 2902
rect 10064 2847 10268 2859
rect 8828 2792 9048 2847
rect 10088 2798 10268 2847
rect 8828 2782 8842 2792
rect 8830 2758 8842 2782
rect 9010 2782 9048 2792
rect 9088 2792 9280 2798
rect 9010 2758 9022 2782
rect 8830 2752 9022 2758
rect 9088 2758 9100 2792
rect 9268 2758 9280 2792
rect 9088 2752 9280 2758
rect 9346 2792 9538 2798
rect 9346 2758 9358 2792
rect 9526 2758 9538 2792
rect 9346 2752 9538 2758
rect 9604 2792 9796 2798
rect 9604 2758 9616 2792
rect 9784 2758 9796 2792
rect 9604 2752 9796 2758
rect 9862 2792 10054 2798
rect 9862 2758 9874 2792
rect 10042 2758 10054 2792
rect 10088 2792 10312 2798
rect 10088 2762 10132 2792
rect 9862 2752 10054 2758
rect 10120 2758 10132 2762
rect 10300 2758 10312 2792
rect 10120 2752 10312 2758
rect 8096 2682 8220 2688
rect 8096 2602 8108 2682
rect 8208 2602 8220 2682
rect 8096 2596 8220 2602
rect 9516 2682 9640 2688
rect 9516 2602 9528 2682
rect 9628 2602 9640 2682
rect 9516 2596 9640 2602
rect 6584 2311 6608 2542
rect 6544 2299 6608 2311
rect 6548 2242 6608 2299
rect 11028 2311 11034 3122
rect 11068 3202 11074 3799
rect 11286 3765 11292 4682
rect 11326 3765 11332 4682
rect 11802 3842 11808 5253
rect 11286 3753 11332 3765
rect 11528 3799 11808 3842
rect 11528 3662 11550 3799
rect 11544 3202 11550 3662
rect 11068 3122 11550 3202
rect 11068 2462 11074 3122
rect 11068 2311 11088 2462
rect 11028 2262 11088 2311
rect 11544 2311 11550 3122
rect 11584 3765 11808 3799
rect 11842 3765 11848 5253
rect 12020 5240 12040 5400
rect 12200 5240 13720 5400
rect 13840 5240 14300 5400
rect 14440 5240 14480 5400
rect 14540 5340 14566 5734
rect 14560 5337 14566 5340
rect 14604 5340 14732 5734
rect 14604 5337 14610 5340
rect 14560 5325 14610 5337
rect 14726 5337 14732 5340
rect 14770 5337 14776 5734
rect 14726 5325 14776 5337
rect 14892 5740 14942 5746
rect 15058 5740 15108 5746
rect 15224 5740 15274 5746
rect 15390 5740 15440 5746
rect 14892 5734 15120 5740
rect 14892 5337 14898 5734
rect 14936 5340 15064 5734
rect 14936 5337 14942 5340
rect 14892 5325 14942 5337
rect 15058 5337 15064 5340
rect 15102 5340 15120 5734
rect 15220 5734 15440 5740
rect 15220 5340 15230 5734
rect 15102 5337 15108 5340
rect 15058 5325 15108 5337
rect 15224 5337 15230 5340
rect 15268 5340 15396 5734
rect 15268 5337 15274 5340
rect 15224 5325 15274 5337
rect 15390 5337 15396 5340
rect 15434 5337 15440 5734
rect 15390 5325 15440 5337
rect 15556 5740 15606 5746
rect 15722 5740 15772 5746
rect 16034 5740 16084 5746
rect 16200 5740 16250 5746
rect 16366 5740 16416 5746
rect 16532 5740 16582 5746
rect 16698 5740 16748 5746
rect 16864 5740 16914 5746
rect 17030 5740 17080 5746
rect 17196 5740 17246 5746
rect 15556 5734 15780 5740
rect 15556 5337 15562 5734
rect 15600 5340 15728 5734
rect 15600 5337 15606 5340
rect 15556 5325 15606 5337
rect 15722 5337 15728 5340
rect 15766 5340 15780 5734
rect 16034 5734 16260 5740
rect 15766 5337 15772 5340
rect 15722 5325 15772 5337
rect 16034 5337 16040 5734
rect 16078 5340 16206 5734
rect 16078 5337 16084 5340
rect 16034 5325 16084 5337
rect 16200 5337 16206 5340
rect 16244 5340 16260 5734
rect 16366 5734 16600 5740
rect 16244 5337 16250 5340
rect 16200 5325 16250 5337
rect 16366 5337 16372 5734
rect 16410 5340 16538 5734
rect 16410 5337 16416 5340
rect 16366 5325 16416 5337
rect 16532 5337 16538 5340
rect 16576 5340 16600 5734
rect 16698 5734 16920 5740
rect 16576 5337 16582 5340
rect 16532 5325 16582 5337
rect 16698 5337 16704 5734
rect 16742 5340 16870 5734
rect 16742 5337 16748 5340
rect 16698 5325 16748 5337
rect 16864 5337 16870 5340
rect 16908 5340 16920 5734
rect 17030 5734 17260 5740
rect 16908 5337 16914 5340
rect 16864 5325 16914 5337
rect 17030 5337 17036 5734
rect 17074 5340 17202 5734
rect 17074 5337 17080 5340
rect 17030 5325 17080 5337
rect 17196 5337 17202 5340
rect 17240 5340 17260 5734
rect 17310 5700 17320 5880
rect 17500 5700 17540 5880
rect 17340 5680 17540 5700
rect 17340 5520 17460 5680
rect 17340 5440 17360 5520
rect 17460 5440 17470 5520
rect 17240 5337 17246 5340
rect 17196 5325 17246 5337
rect 12020 5220 14480 5240
rect 14500 4403 14620 4420
rect 14500 4340 14566 4403
rect 14300 4320 14566 4340
rect 14300 4160 14320 4320
rect 14460 4160 14566 4320
rect 14300 4140 14566 4160
rect 14500 4006 14566 4140
rect 14604 4006 14620 4403
rect 14726 4403 14776 4415
rect 14726 4400 14732 4403
rect 14500 4000 14620 4006
rect 14720 4006 14732 4400
rect 14770 4400 14776 4403
rect 14892 4403 14942 4415
rect 14892 4400 14898 4403
rect 14770 4006 14898 4400
rect 14936 4006 14942 4403
rect 14720 4000 14942 4006
rect 14560 3994 14610 4000
rect 14726 3994 14776 4000
rect 14892 3994 14942 4000
rect 15058 4403 15108 4415
rect 15058 4006 15064 4403
rect 15102 4400 15108 4403
rect 15224 4403 15274 4415
rect 15224 4400 15230 4403
rect 15102 4006 15230 4400
rect 15268 4400 15274 4403
rect 15390 4403 15440 4415
rect 15390 4400 15396 4403
rect 15268 4006 15280 4400
rect 15058 4000 15280 4006
rect 15380 4006 15396 4400
rect 15434 4400 15440 4403
rect 15556 4403 15606 4415
rect 15556 4400 15562 4403
rect 15434 4006 15562 4400
rect 15600 4006 15606 4403
rect 15380 4000 15606 4006
rect 15058 3994 15108 4000
rect 15224 3994 15274 4000
rect 15390 3994 15440 4000
rect 15556 3994 15606 4000
rect 15722 4403 15772 4415
rect 15722 4006 15728 4403
rect 15766 4400 15772 4403
rect 16034 4403 16084 4415
rect 16034 4400 16040 4403
rect 15766 4380 16040 4400
rect 15766 4020 15860 4380
rect 15940 4020 16040 4380
rect 15766 4006 16040 4020
rect 16078 4006 16084 4403
rect 15722 4000 16084 4006
rect 15722 3994 15772 4000
rect 16034 3994 16084 4000
rect 16200 4403 16250 4415
rect 16200 4006 16206 4403
rect 16244 4400 16250 4403
rect 16366 4403 16416 4415
rect 16366 4400 16372 4403
rect 16244 4006 16372 4400
rect 16410 4400 16416 4403
rect 16532 4403 16582 4415
rect 16410 4006 16440 4400
rect 16200 4000 16440 4006
rect 16532 4006 16538 4403
rect 16576 4400 16582 4403
rect 16698 4403 16748 4415
rect 16698 4400 16704 4403
rect 16576 4006 16704 4400
rect 16742 4400 16748 4403
rect 16864 4403 16914 4415
rect 16864 4400 16870 4403
rect 16742 4006 16760 4400
rect 16532 4000 16760 4006
rect 16860 4006 16870 4400
rect 16908 4400 16914 4403
rect 17030 4403 17080 4415
rect 17030 4400 17036 4403
rect 16908 4006 17036 4400
rect 17074 4006 17080 4403
rect 17196 4403 17246 4415
rect 17196 4040 17202 4403
rect 16860 4000 17080 4006
rect 16200 3994 16250 4000
rect 16366 3994 16416 4000
rect 16532 3994 16582 4000
rect 16698 3994 16748 4000
rect 16864 3994 16914 4000
rect 17030 3994 17080 4000
rect 17180 4006 17202 4040
rect 17240 4040 17246 4403
rect 17240 4006 17260 4040
rect 17180 3960 17260 4006
rect 16760 3940 17260 3960
rect 16760 3880 16780 3940
rect 16860 3880 17260 3940
rect 17170 3800 17180 3820
rect 11584 3753 11848 3765
rect 11584 3662 11828 3753
rect 14570 3700 14580 3800
rect 14680 3720 15860 3800
rect 15940 3720 17180 3800
rect 14680 3700 17180 3720
rect 17300 3700 17310 3820
rect 11584 3202 11590 3662
rect 12028 3240 12228 3262
rect 12028 3202 12040 3240
rect 11584 3122 12040 3202
rect 11584 2462 11590 3122
rect 12028 3080 12040 3122
rect 12200 3080 12228 3240
rect 14590 3180 14600 3580
rect 14660 3180 14670 3580
rect 14776 3566 14826 3578
rect 14610 3169 14616 3180
rect 14654 3169 14660 3180
rect 14610 3157 14660 3169
rect 14776 3169 14782 3566
rect 14820 3560 14826 3566
rect 14942 3566 14992 3578
rect 14942 3560 14948 3566
rect 14820 3180 14948 3560
rect 14820 3169 14826 3180
rect 14776 3157 14826 3169
rect 14942 3169 14948 3180
rect 14986 3169 14992 3566
rect 14942 3157 14992 3169
rect 15108 3566 15158 3578
rect 15108 3169 15114 3566
rect 15152 3560 15158 3566
rect 15274 3566 15324 3578
rect 15274 3560 15280 3566
rect 15152 3180 15280 3560
rect 15152 3169 15158 3180
rect 15108 3157 15158 3169
rect 15274 3169 15280 3180
rect 15318 3169 15324 3566
rect 15274 3157 15324 3169
rect 15440 3566 15490 3578
rect 15440 3169 15446 3566
rect 15484 3560 15490 3566
rect 15606 3566 15656 3578
rect 15606 3560 15612 3566
rect 15484 3180 15612 3560
rect 15484 3169 15490 3180
rect 15440 3157 15490 3169
rect 15606 3169 15612 3180
rect 15650 3169 15656 3566
rect 15606 3157 15656 3169
rect 15772 3566 15822 3578
rect 15772 3169 15778 3566
rect 15816 3460 15822 3566
rect 15816 3440 16540 3460
rect 15816 3220 16440 3440
rect 16540 3220 16550 3440
rect 15816 3169 15822 3220
rect 15772 3157 15822 3169
rect 12028 3062 12228 3080
rect 14610 2735 14660 2747
rect 11584 2311 11608 2462
rect 14610 2338 14616 2735
rect 14654 2720 14660 2735
rect 14776 2735 14826 2747
rect 14776 2720 14782 2735
rect 14654 2340 14782 2720
rect 14654 2338 14660 2340
rect 14610 2326 14660 2338
rect 14776 2338 14782 2340
rect 14820 2338 14826 2735
rect 14776 2326 14826 2338
rect 14942 2735 14992 2747
rect 14942 2338 14948 2735
rect 14986 2720 14992 2735
rect 15108 2735 15158 2747
rect 15108 2720 15114 2735
rect 14986 2340 15114 2720
rect 14986 2338 14992 2340
rect 14942 2326 14992 2338
rect 15108 2338 15114 2340
rect 15152 2338 15158 2735
rect 15108 2326 15158 2338
rect 15274 2735 15324 2747
rect 15274 2338 15280 2735
rect 15318 2720 15324 2735
rect 15440 2735 15490 2747
rect 15440 2720 15446 2735
rect 15318 2340 15446 2720
rect 15318 2338 15324 2340
rect 15274 2326 15324 2338
rect 15440 2338 15446 2340
rect 15484 2338 15490 2735
rect 15440 2326 15490 2338
rect 15606 2735 15656 2747
rect 15606 2338 15612 2735
rect 15650 2720 15656 2735
rect 15772 2735 15822 2747
rect 15772 2720 15778 2735
rect 15650 2340 15778 2720
rect 15650 2338 15656 2340
rect 15606 2326 15656 2338
rect 15772 2338 15778 2340
rect 15816 2338 15822 2735
rect 23760 2680 23980 2700
rect 23760 2640 23780 2680
rect 16430 2540 16440 2640
rect 16560 2540 17180 2640
rect 16440 2520 17180 2540
rect 17260 2520 23780 2640
rect 23760 2500 23780 2520
rect 23960 2640 23980 2680
rect 23960 2520 24430 2640
rect 23960 2500 23980 2520
rect 23760 2480 23980 2500
rect 15772 2326 15822 2338
rect 11544 2299 11608 2311
rect 11548 2262 11608 2299
rect 5828 2241 6788 2242
rect 10808 2241 11788 2262
rect 5826 2235 6792 2241
rect 5826 2201 5838 2235
rect 6006 2202 6612 2235
rect 6006 2201 6018 2202
rect 5826 2195 6018 2201
rect 6600 2201 6612 2202
rect 6780 2201 6792 2235
rect 10808 2235 11792 2241
rect 10808 2202 10838 2235
rect 6600 2195 6792 2201
rect 10826 2201 10838 2202
rect 11006 2202 11612 2235
rect 11006 2201 11018 2202
rect 10826 2195 11018 2201
rect 11600 2201 11612 2202
rect 11780 2201 11792 2235
rect 11600 2195 11792 2201
rect 2690 2080 2700 2160
rect 2760 2080 2920 2160
rect 3000 2080 3010 2160
rect 5368 2120 5568 2142
rect 160 1944 480 1970
rect 2670 1960 2680 1980
rect 160 1910 234 1944
rect 402 1910 480 1944
rect 600 1944 2680 1960
rect 600 1920 614 1944
rect 160 1860 480 1910
rect 602 1910 614 1920
rect 782 1920 994 1944
rect 782 1910 794 1920
rect 602 1904 794 1910
rect 982 1910 994 1920
rect 1162 1920 1374 1944
rect 1162 1910 1174 1920
rect 982 1904 1174 1910
rect 1362 1910 1374 1920
rect 1542 1920 1754 1944
rect 1542 1910 1554 1920
rect 1362 1904 1554 1910
rect 1742 1910 1754 1920
rect 1922 1920 2134 1944
rect 1922 1910 1934 1920
rect 1742 1904 1934 1910
rect 2122 1910 2134 1920
rect 2302 1920 2514 1944
rect 2760 1920 2770 1980
rect 5368 1960 5380 2120
rect 5540 2102 5568 2120
rect 5540 2022 7048 2102
rect 7108 2022 7118 2102
rect 5540 1960 5568 2022
rect 2882 1944 3140 1950
rect 2882 1940 2894 1944
rect 2302 1910 2314 1920
rect 2122 1904 2314 1910
rect 2502 1910 2514 1920
rect 2682 1910 2694 1920
rect 2502 1904 2694 1910
rect 2860 1910 2894 1940
rect 3062 1910 3140 1944
rect 5368 1942 5568 1960
rect 2860 1900 3140 1910
rect 546 1870 592 1872
rect 804 1870 850 1872
rect 926 1870 972 1872
rect 1184 1870 1230 1872
rect 160 1684 172 1860
rect 206 1684 430 1860
rect 464 1684 480 1860
rect 530 1690 540 1870
rect 600 1690 610 1870
rect 804 1860 820 1870
rect 960 1860 972 1870
rect 160 1634 480 1684
rect 546 1684 552 1690
rect 586 1684 592 1690
rect 546 1672 592 1684
rect 804 1684 810 1860
rect 966 1684 972 1860
rect 1170 1690 1180 1870
rect 1240 1690 1250 1870
rect 1306 1860 1352 1872
rect 1306 1850 1312 1860
rect 1346 1850 1352 1860
rect 1564 1870 1610 1872
rect 1686 1870 1732 1872
rect 1564 1860 1732 1870
rect 1944 1860 1990 1872
rect 2066 1870 2112 1872
rect 2324 1870 2370 1872
rect 2446 1870 2492 1872
rect 1290 1690 1300 1850
rect 1360 1690 1370 1850
rect 804 1672 820 1684
rect 810 1670 820 1672
rect 960 1672 972 1684
rect 1184 1684 1190 1690
rect 1224 1684 1230 1690
rect 1184 1672 1230 1684
rect 1306 1684 1312 1690
rect 1346 1684 1352 1690
rect 1306 1672 1352 1684
rect 1564 1684 1570 1860
rect 1604 1830 1692 1860
rect 1680 1690 1692 1830
rect 1604 1684 1692 1690
rect 1726 1684 1732 1860
rect 1564 1672 1732 1684
rect 1910 1680 1920 1860
rect 1984 1684 1990 1860
rect 1980 1680 1990 1684
rect 1944 1672 1990 1680
rect 960 1670 970 1672
rect 1580 1670 1720 1672
rect 2030 1670 2040 1870
rect 2120 1670 2130 1870
rect 2324 1860 2492 1870
rect 2324 1684 2330 1860
rect 2364 1850 2452 1860
rect 2364 1684 2370 1690
rect 2324 1672 2370 1684
rect 2446 1684 2452 1690
rect 2486 1684 2492 1860
rect 2704 1860 2750 1872
rect 2704 1850 2710 1860
rect 2446 1672 2492 1684
rect 2670 1670 2680 1850
rect 2744 1684 2750 1860
rect 2740 1670 2750 1684
rect 2820 1860 3140 1900
rect 2820 1684 2832 1860
rect 2866 1684 3090 1860
rect 3124 1684 3140 1860
rect 5368 1820 5568 1822
rect 160 1600 234 1634
rect 402 1600 480 1634
rect 160 1526 480 1600
rect 602 1634 794 1640
rect 602 1600 614 1634
rect 782 1600 794 1634
rect 602 1594 794 1600
rect 982 1634 1174 1640
rect 982 1600 994 1634
rect 1162 1600 1174 1634
rect 982 1594 1174 1600
rect 1362 1634 1554 1640
rect 1362 1600 1374 1634
rect 1542 1600 1554 1634
rect 1362 1594 1554 1600
rect 1742 1634 1934 1640
rect 1742 1600 1754 1634
rect 1922 1600 1934 1634
rect 1742 1594 1934 1600
rect 2122 1634 2314 1640
rect 2122 1600 2134 1634
rect 2302 1600 2314 1634
rect 2122 1594 2314 1600
rect 2502 1634 2694 1640
rect 2502 1600 2514 1634
rect 2682 1600 2694 1634
rect 2502 1594 2694 1600
rect 2820 1634 3140 1684
rect 2820 1600 2894 1634
rect 3062 1600 3140 1634
rect 4980 1800 5568 1820
rect 17170 1800 17180 1860
rect 17240 1840 17250 1860
rect 17240 1834 17260 1840
rect 17242 1800 17260 1834
rect 4980 1640 5000 1800
rect 5120 1782 5568 1800
rect 17196 1794 17254 1800
rect 5120 1662 7908 1782
rect 7988 1662 7998 1782
rect 5120 1640 5568 1662
rect 4980 1622 5568 1640
rect 4980 1620 5560 1622
rect 660 1532 760 1594
rect 1020 1532 1120 1594
rect 1400 1532 1500 1594
rect 1800 1532 1900 1594
rect 2180 1532 2280 1594
rect 2540 1532 2640 1594
rect 160 1492 234 1526
rect 402 1492 480 1526
rect 160 1442 480 1492
rect 602 1526 794 1532
rect 602 1492 614 1526
rect 782 1492 794 1526
rect 602 1486 794 1492
rect 982 1526 1174 1532
rect 982 1492 994 1526
rect 1162 1492 1174 1526
rect 982 1486 1174 1492
rect 1362 1526 1554 1532
rect 1362 1492 1374 1526
rect 1542 1492 1554 1526
rect 1362 1486 1554 1492
rect 1742 1526 1934 1532
rect 1742 1492 1754 1526
rect 1922 1492 1934 1526
rect 1742 1486 1934 1492
rect 2122 1526 2314 1532
rect 2122 1492 2134 1526
rect 2302 1492 2314 1526
rect 2122 1486 2314 1492
rect 2502 1526 2694 1532
rect 2502 1492 2514 1526
rect 2682 1492 2694 1526
rect 2502 1486 2694 1492
rect 2820 1526 3140 1600
rect 12870 1580 12880 1780
rect 13080 1580 14020 1780
rect 14160 1710 14500 1780
rect 14160 1600 16900 1710
rect 16970 1600 16980 1710
rect 14160 1580 14500 1600
rect 14300 1560 14500 1580
rect 2820 1492 2894 1526
rect 3062 1492 3140 1526
rect 1020 1480 1120 1486
rect 1400 1480 1500 1486
rect 1800 1480 1900 1486
rect 2180 1480 2280 1486
rect 2540 1480 2640 1486
rect 546 1450 592 1454
rect 804 1450 850 1454
rect 926 1450 972 1454
rect 1184 1450 1230 1454
rect 160 1266 172 1442
rect 206 1266 430 1442
rect 464 1266 480 1442
rect 160 1216 480 1266
rect 530 1250 540 1450
rect 600 1250 610 1450
rect 804 1442 820 1450
rect 960 1442 972 1450
rect 804 1266 810 1442
rect 966 1266 972 1442
rect 1170 1270 1180 1450
rect 1240 1270 1250 1450
rect 1306 1442 1352 1454
rect 1306 1430 1312 1442
rect 1346 1430 1352 1442
rect 1564 1450 1610 1454
rect 1686 1450 1732 1454
rect 1564 1442 1732 1450
rect 1290 1270 1300 1430
rect 1360 1270 1370 1430
rect 804 1254 820 1266
rect 810 1250 820 1254
rect 960 1254 972 1266
rect 1184 1266 1190 1270
rect 1224 1266 1230 1270
rect 1184 1254 1230 1266
rect 1306 1266 1312 1270
rect 1346 1266 1352 1270
rect 1306 1254 1352 1266
rect 1564 1266 1570 1442
rect 1604 1410 1692 1442
rect 1604 1266 1692 1270
rect 1726 1266 1732 1442
rect 1944 1442 1990 1454
rect 2066 1450 2112 1454
rect 2324 1450 2370 1454
rect 2446 1450 2492 1454
rect 2704 1450 2750 1454
rect 1944 1440 1950 1442
rect 1564 1254 1732 1266
rect 1910 1260 1920 1440
rect 1984 1266 1990 1442
rect 1980 1260 1990 1266
rect 1944 1254 1990 1260
rect 960 1250 970 1254
rect 1580 1250 1720 1254
rect 2050 1250 2060 1450
rect 2140 1250 2150 1450
rect 2324 1442 2492 1450
rect 2324 1266 2330 1442
rect 2364 1430 2452 1442
rect 2364 1266 2370 1270
rect 2324 1254 2370 1266
rect 2446 1266 2452 1270
rect 2486 1266 2492 1442
rect 2690 1270 2700 1450
rect 2760 1270 2770 1450
rect 2820 1442 3140 1492
rect 2446 1254 2492 1266
rect 2704 1266 2710 1270
rect 2744 1266 2750 1270
rect 2704 1254 2750 1266
rect 2820 1266 2832 1442
rect 2866 1266 3090 1442
rect 3124 1266 3140 1442
rect 160 1182 234 1216
rect 402 1182 480 1216
rect 160 1108 480 1182
rect 602 1216 794 1222
rect 602 1182 614 1216
rect 782 1182 794 1216
rect 602 1176 794 1182
rect 982 1216 1174 1222
rect 982 1182 994 1216
rect 1162 1182 1174 1216
rect 982 1176 1174 1182
rect 1362 1216 1554 1222
rect 1362 1182 1374 1216
rect 1542 1182 1554 1216
rect 1362 1176 1554 1182
rect 1742 1216 1934 1222
rect 1742 1182 1754 1216
rect 1922 1182 1934 1216
rect 1742 1176 1934 1182
rect 2122 1216 2314 1222
rect 2122 1182 2134 1216
rect 2302 1182 2314 1216
rect 2122 1176 2314 1182
rect 2502 1216 2694 1222
rect 2502 1182 2514 1216
rect 2682 1182 2694 1216
rect 2502 1176 2694 1182
rect 2820 1216 3140 1266
rect 14300 1420 14500 1460
rect 14300 1280 14340 1420
rect 14460 1400 14500 1420
rect 14460 1369 16714 1400
rect 14460 1335 14627 1369
rect 14661 1335 14719 1369
rect 14753 1335 14811 1369
rect 14845 1335 14903 1369
rect 14937 1335 14995 1369
rect 15029 1335 15087 1369
rect 15121 1335 15179 1369
rect 15213 1335 15271 1369
rect 15305 1335 15363 1369
rect 15397 1335 15455 1369
rect 15489 1335 15547 1369
rect 15581 1335 15639 1369
rect 15673 1335 15731 1369
rect 15765 1335 15823 1369
rect 15857 1335 15915 1369
rect 15949 1335 16007 1369
rect 16041 1335 16099 1369
rect 16133 1335 16191 1369
rect 16225 1335 16283 1369
rect 16317 1335 16375 1369
rect 16409 1335 16467 1369
rect 16501 1335 16559 1369
rect 16593 1335 16651 1369
rect 16685 1335 16714 1369
rect 14460 1304 16714 1335
rect 14460 1300 14640 1304
rect 14300 1260 14430 1280
rect 14420 1250 14430 1260
rect 14500 1250 14520 1300
rect 14420 1220 14520 1250
rect 2820 1182 2894 1216
rect 3062 1182 3140 1216
rect 660 1114 760 1176
rect 1020 1114 1120 1176
rect 1400 1114 1500 1176
rect 1800 1114 1900 1176
rect 2180 1114 2280 1176
rect 2540 1114 2640 1176
rect 160 1074 234 1108
rect 402 1074 480 1108
rect 160 1024 480 1074
rect 602 1108 794 1114
rect 602 1074 614 1108
rect 782 1074 794 1108
rect 602 1068 794 1074
rect 982 1108 1174 1114
rect 982 1074 994 1108
rect 1162 1074 1174 1108
rect 982 1068 1174 1074
rect 1362 1108 1554 1114
rect 1362 1074 1374 1108
rect 1542 1074 1554 1108
rect 1362 1068 1554 1074
rect 1742 1108 1934 1114
rect 1742 1074 1754 1108
rect 1922 1074 1934 1108
rect 1742 1068 1934 1074
rect 2122 1108 2314 1114
rect 2122 1074 2134 1108
rect 2302 1074 2314 1108
rect 2122 1068 2314 1074
rect 2502 1108 2694 1114
rect 2502 1074 2514 1108
rect 2682 1074 2694 1108
rect 2502 1068 2694 1074
rect 2820 1108 3140 1182
rect 14789 1199 14847 1205
rect 14789 1165 14801 1199
rect 14835 1196 14847 1199
rect 15167 1199 15225 1205
rect 15167 1196 15179 1199
rect 14835 1168 15179 1196
rect 14835 1165 14847 1168
rect 14789 1159 14847 1165
rect 15167 1165 15179 1168
rect 15213 1196 15225 1199
rect 15791 1199 15849 1205
rect 15791 1196 15803 1199
rect 15213 1168 15803 1196
rect 15213 1165 15225 1168
rect 15167 1159 15225 1165
rect 15791 1165 15803 1168
rect 15837 1165 15849 1199
rect 17070 1180 17080 1760
rect 17140 1753 17180 1760
rect 17140 1741 17204 1753
rect 17140 1180 17164 1741
rect 15791 1159 15849 1165
rect 17158 1165 17164 1180
rect 17198 1165 17204 1741
rect 17158 1153 17204 1165
rect 17246 1741 17292 1753
rect 17246 1165 17252 1741
rect 17286 1740 17292 1741
rect 17354 1740 17406 1752
rect 17286 1180 17360 1740
rect 17400 1720 17440 1740
rect 17440 1640 17450 1720
rect 17400 1600 17440 1640
rect 17440 1520 17450 1600
rect 17400 1460 17440 1520
rect 17440 1380 17450 1460
rect 17400 1320 17440 1380
rect 17440 1240 17450 1320
rect 17400 1180 17440 1240
rect 17286 1165 17292 1180
rect 17354 1168 17406 1180
rect 17246 1153 17292 1165
rect 2820 1074 2894 1108
rect 3062 1074 3140 1108
rect 13080 1100 14500 1120
rect 17196 1106 17254 1112
rect 17196 1100 17208 1106
rect 17242 1100 17254 1106
rect 546 1030 592 1036
rect 804 1030 850 1036
rect 926 1030 972 1036
rect 1184 1030 1230 1036
rect 160 848 172 1024
rect 206 848 430 1024
rect 464 848 480 1024
rect 530 850 540 1030
rect 600 850 610 1030
rect 804 1024 820 1030
rect 960 1024 972 1030
rect 160 798 480 848
rect 546 848 552 850
rect 586 848 592 850
rect 546 836 592 848
rect 804 848 810 1024
rect 966 848 972 1024
rect 1170 850 1180 1030
rect 1240 850 1250 1030
rect 1306 1024 1352 1036
rect 1306 1010 1312 1024
rect 1346 1010 1352 1024
rect 1564 1030 1610 1036
rect 1686 1030 1732 1036
rect 1564 1024 1732 1030
rect 1290 850 1300 1010
rect 1360 850 1370 1010
rect 804 836 820 848
rect 810 830 820 836
rect 960 836 972 848
rect 1184 848 1190 850
rect 1224 848 1230 850
rect 1184 836 1230 848
rect 1306 848 1312 850
rect 1346 848 1352 850
rect 1306 836 1352 848
rect 1564 848 1570 1024
rect 1604 990 1692 1024
rect 1604 848 1692 850
rect 1726 848 1732 1024
rect 1944 1024 1990 1036
rect 2066 1030 2112 1036
rect 2324 1030 2370 1036
rect 2446 1030 2492 1036
rect 2704 1030 2750 1036
rect 1944 1020 1950 1024
rect 1564 836 1732 848
rect 1910 840 1920 1020
rect 1984 848 1990 1024
rect 2050 850 2060 1030
rect 2120 850 2130 1030
rect 2324 1024 2492 1030
rect 1980 840 1990 848
rect 1944 836 1990 840
rect 2066 848 2072 850
rect 2106 848 2112 850
rect 2066 836 2112 848
rect 2324 848 2330 1024
rect 2364 1010 2452 1024
rect 2364 848 2370 850
rect 2324 836 2370 848
rect 2446 848 2452 850
rect 2486 848 2492 1024
rect 2690 850 2700 1030
rect 2760 850 2770 1030
rect 2820 1024 3140 1074
rect 2446 836 2492 848
rect 2704 848 2710 850
rect 2744 848 2750 850
rect 2704 836 2750 848
rect 2820 848 2832 1024
rect 2866 848 3090 1024
rect 3124 848 3140 1024
rect 13070 920 13080 1100
rect 13260 1080 14500 1100
rect 14614 1080 14666 1092
rect 13260 1020 14620 1080
rect 14660 1020 14666 1080
rect 14708 1063 14766 1069
rect 14708 1029 14720 1063
rect 14754 1060 14766 1063
rect 15075 1063 15133 1069
rect 15075 1060 15087 1063
rect 14754 1032 15087 1060
rect 14754 1029 14766 1032
rect 14708 1023 14766 1029
rect 15075 1029 15087 1032
rect 15121 1060 15133 1063
rect 15791 1063 15849 1069
rect 15791 1060 15803 1063
rect 15121 1032 15803 1060
rect 15121 1029 15133 1032
rect 15075 1023 15133 1029
rect 15791 1029 15803 1032
rect 15837 1029 15849 1063
rect 15791 1023 15849 1029
rect 16007 1058 16065 1064
rect 16007 1024 16019 1058
rect 16053 1024 16065 1058
rect 13260 920 14500 1020
rect 14614 1008 14666 1020
rect 16007 1001 16065 1024
rect 16638 1060 16702 1066
rect 16890 1060 16900 1080
rect 16638 1020 16650 1060
rect 16690 1020 16900 1060
rect 16638 1014 16702 1020
rect 15347 1000 15477 1001
rect 14880 930 14890 1000
rect 14970 930 14980 1000
rect 15330 940 15340 1000
rect 15400 995 15477 1000
rect 15400 961 15431 995
rect 15465 992 15477 995
rect 16007 995 16125 1001
rect 16890 1000 16900 1020
rect 16980 1000 16990 1080
rect 17180 1060 17200 1100
rect 17190 1040 17200 1060
rect 17260 1040 17270 1100
rect 16007 992 16079 995
rect 15465 964 16079 992
rect 15465 961 15477 964
rect 15400 955 15477 961
rect 16067 961 16079 964
rect 16113 961 16125 995
rect 16067 955 16125 961
rect 16328 960 16412 966
rect 15400 940 15410 955
rect 16328 900 16340 960
rect 16400 900 16780 960
rect 16860 900 16870 960
rect 16328 894 16412 900
rect 960 830 970 836
rect 1580 830 1720 836
rect 160 764 234 798
rect 402 764 480 798
rect 160 690 480 764
rect 602 798 794 804
rect 602 764 614 798
rect 782 764 794 798
rect 602 758 794 764
rect 982 798 1174 804
rect 982 764 994 798
rect 1162 764 1174 798
rect 982 758 1174 764
rect 1362 798 1554 804
rect 1362 764 1374 798
rect 1542 764 1554 798
rect 1362 758 1554 764
rect 1742 798 1934 804
rect 1742 764 1754 798
rect 1922 764 1934 798
rect 1742 758 1934 764
rect 2122 798 2314 804
rect 2122 764 2134 798
rect 2302 764 2314 798
rect 2122 758 2314 764
rect 2502 798 2694 804
rect 2502 764 2514 798
rect 2682 764 2694 798
rect 2502 758 2694 764
rect 2820 798 3140 848
rect 2820 764 2894 798
rect 3062 764 3140 798
rect 660 696 760 758
rect 1020 696 1120 758
rect 1400 696 1500 758
rect 1800 696 1900 758
rect 2180 696 2280 758
rect 2540 696 2640 758
rect 160 656 234 690
rect 402 656 480 690
rect 160 606 480 656
rect 602 690 794 696
rect 602 656 614 690
rect 782 656 794 690
rect 602 650 794 656
rect 982 690 1174 696
rect 982 656 994 690
rect 1162 656 1174 690
rect 982 650 1174 656
rect 1362 690 1554 696
rect 1362 656 1374 690
rect 1542 656 1554 690
rect 1362 650 1554 656
rect 1742 690 1934 696
rect 1742 656 1754 690
rect 1922 656 1934 690
rect 1742 650 1934 656
rect 2122 690 2314 696
rect 2122 656 2134 690
rect 2302 656 2314 690
rect 2122 650 2314 656
rect 2502 690 2694 696
rect 2502 656 2514 690
rect 2682 656 2694 690
rect 2502 650 2694 656
rect 2820 690 3140 764
rect 14598 840 16714 856
rect 14598 760 14620 840
rect 14700 825 16714 840
rect 14700 791 14719 825
rect 14753 791 14811 825
rect 14845 791 14903 825
rect 14937 791 14995 825
rect 15029 791 15087 825
rect 15121 791 15179 825
rect 15213 791 15271 825
rect 15305 791 15363 825
rect 15397 791 15455 825
rect 15489 791 15547 825
rect 15581 791 15639 825
rect 15673 791 15731 825
rect 15765 791 15823 825
rect 15857 791 15915 825
rect 15949 791 16007 825
rect 16041 791 16099 825
rect 16133 791 16191 825
rect 16225 791 16283 825
rect 16317 791 16375 825
rect 16409 791 16467 825
rect 16501 791 16559 825
rect 16593 791 16651 825
rect 16685 791 16714 825
rect 14700 760 16714 791
rect 17190 760 17200 780
rect 17180 720 17200 760
rect 17260 720 17270 780
rect 2820 656 2894 690
rect 3062 656 3140 690
rect 14890 660 14900 720
rect 14960 710 17130 720
rect 14960 660 17060 710
rect 546 610 592 618
rect 804 610 850 618
rect 926 610 972 618
rect 1184 610 1230 618
rect 160 430 172 606
rect 206 430 430 606
rect 464 430 480 606
rect 530 430 540 610
rect 600 430 610 610
rect 804 606 820 610
rect 960 606 972 610
rect 804 430 810 606
rect 966 430 972 606
rect 1170 430 1180 610
rect 1240 430 1250 610
rect 1306 606 1352 618
rect 1306 590 1312 606
rect 1346 590 1352 606
rect 1564 610 1610 618
rect 1686 610 1732 618
rect 1564 606 1732 610
rect 1290 430 1300 590
rect 1360 430 1370 590
rect 1564 430 1570 606
rect 1604 570 1692 606
rect 1726 430 1732 606
rect 1944 606 1990 618
rect 2066 610 2112 618
rect 2324 610 2370 618
rect 2446 610 2492 618
rect 2704 610 2750 618
rect 1944 600 1950 606
rect 160 380 480 430
rect 546 418 592 430
rect 804 418 850 430
rect 926 418 972 430
rect 1184 418 1230 430
rect 1306 418 1352 430
rect 1564 418 1732 430
rect 1910 420 1920 600
rect 1984 430 1990 606
rect 2050 430 2060 610
rect 2120 430 2130 610
rect 2324 606 2492 610
rect 2324 430 2330 606
rect 2364 590 2452 606
rect 2486 430 2492 606
rect 2690 430 2700 610
rect 2760 430 2770 610
rect 2820 606 3140 656
rect 17050 650 17060 660
rect 17120 660 17130 710
rect 17196 712 17208 720
rect 17242 712 17254 720
rect 17196 706 17254 712
rect 17158 662 17204 674
rect 17158 660 17164 662
rect 17120 650 17164 660
rect 2820 430 2832 606
rect 2866 430 3090 606
rect 3124 430 3140 606
rect 1980 420 1990 430
rect 1944 418 1990 420
rect 2066 418 2112 430
rect 2324 418 2370 430
rect 2446 418 2492 430
rect 2704 418 2750 430
rect 1580 410 1720 418
rect 160 346 234 380
rect 402 346 480 380
rect 160 240 480 346
rect 602 380 794 386
rect 602 346 614 380
rect 782 346 794 380
rect 602 340 794 346
rect 982 380 1174 386
rect 982 346 994 380
rect 1162 346 1174 380
rect 982 340 1174 346
rect 1362 380 1554 386
rect 1362 346 1374 380
rect 1542 346 1554 380
rect 1362 340 1554 346
rect 1742 380 1934 386
rect 1742 346 1754 380
rect 1922 346 1934 380
rect 1742 340 1934 346
rect 2122 380 2314 386
rect 2122 346 2134 380
rect 2302 346 2314 380
rect 2122 340 2314 346
rect 2502 380 2694 386
rect 2502 346 2514 380
rect 2682 346 2694 380
rect 2502 340 2694 346
rect 2820 380 3140 430
rect 2820 346 2894 380
rect 3062 346 3140 380
rect 14300 540 14500 560
rect 14300 360 14340 540
rect 14460 500 14500 540
rect 14460 440 15340 500
rect 15400 440 15410 500
rect 17070 486 17164 650
rect 17198 486 17204 662
rect 17070 480 17204 486
rect 17158 474 17204 480
rect 17246 662 17292 674
rect 17246 486 17252 662
rect 17286 660 17292 662
rect 17286 640 17460 660
rect 17286 620 17360 640
rect 17400 620 17460 640
rect 17286 486 17320 620
rect 17246 480 17320 486
rect 17420 480 17460 620
rect 17246 474 17292 480
rect 17340 460 17460 480
rect 17196 440 17254 442
rect 14460 360 14500 440
rect 17180 436 17260 440
rect 17180 402 17208 436
rect 17242 402 17260 436
rect 17180 400 17260 402
rect 17196 396 17254 400
rect 160 200 220 240
rect 440 210 480 240
rect 1088 240 1332 246
rect 1088 210 1100 240
rect 440 200 1100 210
rect 1320 210 1332 240
rect 2008 240 2252 246
rect 2008 210 2020 240
rect 1320 200 1580 210
rect 160 190 1580 200
rect 160 160 840 190
rect 160 40 200 160
rect 480 90 840 160
rect 940 90 1580 190
rect 480 70 1580 90
rect 1700 200 2020 210
rect 2240 210 2252 240
rect 2820 240 3140 346
rect 2820 210 2860 240
rect 2240 200 2340 210
rect 1700 70 2340 200
rect 2480 200 2860 210
rect 3080 200 3140 240
rect 2480 70 3140 200
rect 15720 160 15920 200
rect 480 40 3140 70
rect 160 0 3140 40
rect 14580 20 14600 160
rect 14700 140 17420 160
rect 14700 20 15640 140
rect 15900 20 17320 140
rect 17420 20 17430 140
rect 14580 0 17420 20
rect 16030 -20 16190 0
rect 58 -1616 16098 -1596
rect 58 -1756 198 -1616
rect -62 -1916 198 -1756
rect 458 -1636 16098 -1616
rect 458 -1658 15678 -1636
rect 458 -1718 8128 -1658
rect 8188 -1718 9548 -1658
rect 9608 -1718 15678 -1658
rect 458 -1876 15678 -1718
rect 15878 -1876 16098 -1636
rect 458 -1916 16098 -1876
rect -62 -1956 16098 -1916
rect 58 -2036 16098 -1956
rect 4958 -2160 5158 -2156
rect 4358 -2196 4558 -2176
rect 4348 -2296 4358 -2196
rect 4558 -2296 4568 -2196
rect 4360 -2580 4560 -2296
rect 4950 -2300 4960 -2160
rect 5160 -2300 5170 -2160
rect 13078 -2176 13278 -2156
rect 14298 -2176 14498 -2156
rect 13078 -2276 13098 -2176
rect 13258 -2276 13278 -2176
rect 4958 -2576 5158 -2300
rect 13078 -2576 13278 -2276
rect 13698 -2196 13858 -2176
rect 13698 -2276 13718 -2196
rect 13838 -2276 13858 -2196
rect 13698 -2376 13858 -2276
rect 14008 -2296 14018 -2176
rect 14178 -2296 14188 -2176
rect 14298 -2276 14318 -2176
rect 14478 -2276 14498 -2176
rect 13658 -2576 13858 -2376
rect 14018 -2376 14178 -2296
rect 14298 -2376 14498 -2276
rect 14018 -2576 14218 -2376
rect 14278 -2576 14478 -2376
<< via1 >>
rect 6940 6880 7260 7160
rect 12880 6560 13080 6760
rect 320 5300 400 5400
rect 1600 5300 1720 5400
rect 3500 5320 4000 5480
rect 6288 5442 6348 5562
rect 8188 5442 8288 5542
rect 8760 5540 8960 5900
rect 9328 5442 9428 5542
rect 11268 5422 11328 5522
rect 4040 5300 4140 5400
rect 1600 4840 1720 4960
rect 2360 4592 2406 4800
rect 2406 4592 2440 4800
rect 2360 4580 2440 4592
rect 3280 4620 3380 4740
rect 4040 4840 4140 4960
rect 2620 4533 2720 4540
rect 2620 4499 2720 4533
rect 2620 4480 2720 4499
rect 320 4271 400 4300
rect 320 4220 388 4271
rect 388 4220 400 4271
rect 2360 4200 2440 4300
rect 2920 4180 3020 4280
rect 840 3853 940 3860
rect 840 3819 940 3853
rect 840 3800 940 3819
rect 2620 3853 2720 3860
rect 2620 3819 2630 3853
rect 2630 3819 2720 3853
rect 2620 3800 2720 3819
rect 6268 4882 6292 5122
rect 6292 4882 6326 5122
rect 6326 4882 6368 5122
rect 2620 3420 2720 3540
rect 2620 2613 2700 2780
rect 3280 2940 3360 3040
rect 3360 2940 3400 3040
rect 4380 2900 4560 3100
rect 5380 2920 5540 3080
rect 2620 2580 2700 2613
rect 2040 2420 2100 2480
rect 2920 2420 3020 2480
rect 540 2240 600 2320
rect 840 2240 940 2300
rect 1180 2240 1240 2320
rect 1300 2280 1360 2360
rect 1940 2280 2000 2360
rect 2620 2280 2720 2360
rect 8188 5253 8288 5282
rect 8188 5202 8226 5253
rect 8226 5202 8260 5253
rect 8260 5202 8288 5253
rect 8468 5111 8484 5182
rect 8484 5111 8518 5182
rect 8518 5111 8548 5182
rect 8468 5082 8548 5111
rect 9108 5165 9114 5242
rect 9114 5165 9148 5242
rect 9148 5165 9188 5242
rect 9108 5162 9188 5165
rect 9348 5199 9428 5202
rect 9348 5111 9372 5199
rect 9372 5111 9406 5199
rect 9406 5111 9428 5199
rect 9348 5082 9428 5111
rect 8768 4742 8848 4822
rect 10528 4742 10608 4822
rect 8768 4682 8848 4702
rect 8768 4648 8784 4682
rect 8784 4648 8818 4682
rect 8818 4648 8848 4682
rect 8768 4642 8848 4648
rect 8468 4522 8548 4602
rect 9108 4522 9188 4602
rect 8808 4339 8832 4402
rect 8832 4339 8866 4402
rect 8866 4339 8868 4402
rect 8808 4322 8868 4339
rect 9108 4222 9168 4282
rect 7048 4102 7108 4162
rect 9108 4102 9168 4162
rect 8388 4002 8468 4062
rect 8808 4002 8868 4062
rect 7908 3773 7912 3822
rect 7912 3773 7988 3822
rect 7908 3742 7988 3773
rect 8108 3719 8136 3802
rect 8136 3719 8170 3802
rect 8170 3719 8208 3802
rect 8108 3702 8208 3719
rect 8388 3861 8448 3862
rect 8388 3773 8394 3861
rect 8394 3773 8428 3861
rect 8428 3773 8448 3861
rect 8388 3762 8448 3773
rect 8868 3622 8928 3682
rect 9148 3622 9208 3802
rect 8868 3062 8928 3122
rect 10188 3502 10248 3562
rect 9528 2862 9554 3102
rect 9554 2862 9588 3102
rect 11268 4682 11292 5242
rect 11292 4682 11326 5242
rect 11326 4682 11328 5242
rect 10208 3122 10268 3182
rect 10528 3142 10588 3202
rect 8108 2602 8208 2682
rect 9528 2602 9628 2682
rect 12040 5240 12200 5400
rect 13720 5240 13840 5400
rect 14300 5240 14440 5400
rect 17320 5700 17500 5880
rect 17360 5440 17460 5520
rect 14320 4160 14460 4320
rect 15860 4020 15940 4380
rect 16780 3880 16860 3940
rect 14580 3700 14680 3800
rect 15860 3720 15940 3800
rect 17180 3700 17300 3820
rect 12040 3080 12200 3240
rect 14600 3566 14660 3580
rect 14600 3180 14616 3566
rect 14616 3180 14654 3566
rect 14654 3180 14660 3566
rect 16440 3220 16540 3440
rect 16440 2540 16560 2640
rect 17180 2520 17260 2640
rect 23780 2500 23960 2680
rect 2700 2080 2760 2160
rect 2920 2080 3000 2160
rect 2680 1944 2760 1980
rect 2680 1920 2682 1944
rect 2682 1920 2760 1944
rect 5380 1960 5540 2120
rect 7048 2022 7108 2102
rect 540 1860 600 1870
rect 540 1690 552 1860
rect 552 1690 586 1860
rect 586 1690 600 1860
rect 820 1860 960 1870
rect 820 1684 844 1860
rect 844 1684 932 1860
rect 932 1684 960 1860
rect 1180 1860 1240 1870
rect 1180 1690 1190 1860
rect 1190 1690 1224 1860
rect 1224 1690 1240 1860
rect 1300 1690 1312 1850
rect 1312 1690 1346 1850
rect 1346 1690 1360 1850
rect 820 1670 960 1684
rect 1580 1690 1604 1830
rect 1604 1690 1680 1830
rect 1920 1684 1950 1860
rect 1950 1684 1980 1860
rect 1920 1680 1980 1684
rect 2040 1860 2120 1870
rect 2040 1684 2072 1860
rect 2072 1684 2106 1860
rect 2106 1684 2120 1860
rect 2040 1670 2120 1684
rect 2340 1690 2364 1850
rect 2364 1690 2452 1850
rect 2452 1690 2460 1850
rect 2680 1684 2710 1850
rect 2710 1684 2740 1850
rect 2680 1670 2740 1684
rect 17180 1834 17240 1860
rect 17180 1800 17208 1834
rect 17208 1800 17240 1834
rect 5000 1640 5120 1800
rect 7908 1662 7988 1782
rect 12880 1580 13080 1780
rect 14020 1580 14160 1780
rect 16900 1600 16970 1710
rect 540 1442 600 1450
rect 540 1266 552 1442
rect 552 1266 586 1442
rect 586 1266 600 1442
rect 540 1250 600 1266
rect 820 1442 960 1450
rect 820 1266 844 1442
rect 844 1266 932 1442
rect 932 1266 960 1442
rect 1180 1442 1240 1450
rect 1180 1270 1190 1442
rect 1190 1270 1224 1442
rect 1224 1270 1240 1442
rect 1300 1270 1312 1430
rect 1312 1270 1346 1430
rect 1346 1270 1360 1430
rect 820 1250 960 1266
rect 1600 1270 1604 1410
rect 1604 1270 1692 1410
rect 1692 1270 1700 1410
rect 1920 1266 1950 1440
rect 1950 1266 1980 1440
rect 1920 1260 1980 1266
rect 2060 1442 2140 1450
rect 2060 1266 2072 1442
rect 2072 1266 2106 1442
rect 2106 1266 2140 1442
rect 2060 1250 2140 1266
rect 2340 1270 2364 1430
rect 2364 1270 2452 1430
rect 2452 1270 2460 1430
rect 2700 1442 2760 1450
rect 2700 1270 2710 1442
rect 2710 1270 2744 1442
rect 2744 1270 2760 1442
rect 14340 1300 14460 1420
rect 14340 1280 14430 1300
rect 14430 1280 14460 1300
rect 17080 1180 17140 1760
rect 17360 1640 17400 1720
rect 17400 1640 17440 1720
rect 17360 1520 17400 1600
rect 17400 1520 17440 1600
rect 17360 1380 17400 1460
rect 17400 1380 17440 1460
rect 17360 1240 17400 1320
rect 17400 1240 17440 1320
rect 540 1024 600 1030
rect 540 850 552 1024
rect 552 850 586 1024
rect 586 850 600 1024
rect 820 1024 960 1030
rect 820 848 844 1024
rect 844 848 932 1024
rect 932 848 960 1024
rect 1180 1024 1240 1030
rect 1180 850 1190 1024
rect 1190 850 1224 1024
rect 1224 850 1240 1024
rect 1300 850 1312 1010
rect 1312 850 1346 1010
rect 1346 850 1360 1010
rect 820 830 960 848
rect 1600 850 1604 990
rect 1604 850 1692 990
rect 1692 850 1700 990
rect 1920 848 1950 1020
rect 1950 848 1980 1020
rect 2060 1024 2120 1030
rect 2060 850 2072 1024
rect 2072 850 2106 1024
rect 2106 850 2120 1024
rect 1920 840 1980 848
rect 2340 850 2364 1010
rect 2364 850 2452 1010
rect 2452 850 2460 1010
rect 2700 1024 2760 1030
rect 2700 850 2710 1024
rect 2710 850 2744 1024
rect 2744 850 2760 1024
rect 13080 920 13260 1100
rect 14890 990 14970 1000
rect 14890 950 14900 990
rect 14900 950 14960 990
rect 14960 950 14970 990
rect 14890 930 14970 950
rect 15340 995 15400 1000
rect 15340 961 15359 995
rect 15359 961 15393 995
rect 15393 961 15400 995
rect 16900 1000 16980 1080
rect 17200 1072 17208 1100
rect 17208 1072 17242 1100
rect 17242 1072 17260 1100
rect 17200 1040 17260 1072
rect 15340 940 15400 961
rect 16780 900 16860 960
rect 14620 825 14700 840
rect 14620 791 14627 825
rect 14627 791 14661 825
rect 14661 791 14700 825
rect 14620 760 14700 791
rect 17200 746 17260 780
rect 17200 720 17208 746
rect 17208 720 17242 746
rect 17242 720 17260 746
rect 14900 660 14960 720
rect 540 606 600 610
rect 540 430 552 606
rect 552 430 586 606
rect 586 430 600 606
rect 820 606 960 610
rect 820 430 844 606
rect 844 430 932 606
rect 932 430 960 606
rect 1180 606 1240 610
rect 1180 430 1190 606
rect 1190 430 1224 606
rect 1224 430 1240 606
rect 1300 430 1312 590
rect 1312 430 1346 590
rect 1346 430 1360 590
rect 1600 430 1604 570
rect 1604 430 1692 570
rect 1692 430 1700 570
rect 1920 430 1950 600
rect 1950 430 1980 600
rect 2060 606 2120 610
rect 2060 430 2072 606
rect 2072 430 2106 606
rect 2106 430 2120 606
rect 2340 430 2364 590
rect 2364 430 2452 590
rect 2452 430 2460 590
rect 2700 606 2760 610
rect 2700 430 2710 606
rect 2710 430 2744 606
rect 2744 430 2760 606
rect 17060 650 17120 710
rect 1920 420 1980 430
rect 14340 360 14460 540
rect 15340 440 15400 500
rect 17320 480 17360 620
rect 17360 480 17400 620
rect 17400 480 17420 620
rect 200 40 480 160
rect 840 90 940 190
rect 1580 70 1700 210
rect 2340 70 2480 210
rect 14600 20 14700 160
rect 15640 20 15900 140
rect 17320 20 17420 140
rect 198 -1916 458 -1616
rect 8128 -1718 8188 -1658
rect 9548 -1718 9608 -1658
rect 15678 -1876 15878 -1636
rect 4358 -2296 4558 -2196
rect 4960 -2300 5160 -2160
rect 13098 -2276 13258 -2176
rect 13718 -2276 13838 -2196
rect 14018 -2296 14178 -2176
rect 14318 -2276 14478 -2176
<< metal2 >>
rect 6940 7160 7260 7170
rect 6940 6870 7260 6880
rect 12880 6760 13100 6780
rect 13080 6560 13100 6760
rect 8760 5900 8960 5910
rect 6288 5562 6348 5572
rect 3500 5480 4000 5490
rect 320 5400 400 5410
rect 320 4300 400 5300
rect 1600 5400 1720 5410
rect 6268 5442 6288 5562
rect 6348 5442 6368 5562
rect 3500 5310 4000 5320
rect 4040 5400 4140 5410
rect 1600 4960 1720 5300
rect 1600 4830 1720 4840
rect 4040 4960 4140 5300
rect 6268 5122 6368 5442
rect 8188 5542 8288 5552
rect 8760 5530 8960 5540
rect 9328 5542 9428 5552
rect 8188 5282 8288 5442
rect 9108 5242 9188 5252
rect 8188 5192 8288 5202
rect 6268 4872 6368 4882
rect 8468 5182 8548 5202
rect 4040 4830 4140 4840
rect 320 4210 400 4220
rect 2360 4800 2440 4810
rect 2360 4300 2440 4580
rect 3280 4740 3400 4760
rect 3380 4620 3400 4740
rect 2360 4190 2440 4200
rect 2620 4540 2720 4550
rect 840 3860 940 3870
rect 540 2320 600 2330
rect 540 1870 600 2240
rect 840 2300 940 3800
rect 2620 3860 2720 4480
rect 2620 3540 2720 3800
rect 2620 2780 2720 3420
rect 2700 2580 2720 2780
rect 2040 2480 2100 2490
rect 1300 2360 1360 2370
rect 840 2230 940 2240
rect 1180 2320 1240 2330
rect 540 1450 600 1690
rect 540 1030 600 1250
rect 540 610 600 850
rect 540 410 600 430
rect 820 1870 960 1880
rect 820 1450 960 1670
rect 820 1030 960 1250
rect 820 610 960 830
rect 820 190 960 430
rect 1180 1870 1240 2240
rect 1180 1450 1240 1690
rect 1180 1030 1240 1270
rect 1180 610 1240 850
rect 1180 410 1240 430
rect 1300 1850 1360 2280
rect 1940 2360 2000 2370
rect 1940 1870 2000 2280
rect 1920 1860 2000 1870
rect 1300 1430 1360 1690
rect 1300 1010 1360 1270
rect 1300 590 1360 850
rect 1300 410 1360 430
rect 1580 1830 1700 1850
rect 1680 1690 1700 1830
rect 1580 1410 1700 1690
rect 1980 1680 2000 1860
rect 1920 1670 2000 1680
rect 1940 1450 2000 1670
rect 1580 1270 1600 1410
rect 1580 990 1700 1270
rect 1920 1440 2000 1450
rect 1980 1260 2000 1440
rect 1920 1250 2000 1260
rect 1940 1030 2000 1250
rect 1580 850 1600 990
rect 1580 570 1700 850
rect 1920 1020 2000 1030
rect 1980 840 2000 1020
rect 1920 830 2000 840
rect 1940 610 2000 830
rect 1580 430 1600 570
rect 160 160 500 180
rect 160 40 200 160
rect 480 40 500 160
rect 820 90 840 190
rect 940 90 960 190
rect 820 70 960 90
rect 1580 210 1700 430
rect 1920 600 2000 610
rect 1980 420 2000 600
rect 1920 410 2000 420
rect 2040 1880 2100 2420
rect 2620 2360 2720 2580
rect 2620 2270 2720 2280
rect 2920 4280 3020 4290
rect 2920 2480 3020 4180
rect 3280 3040 3400 4620
rect 8468 4602 8548 5082
rect 8768 4822 8848 4832
rect 8768 4702 8848 4742
rect 8768 4632 8848 4642
rect 8468 4512 8548 4522
rect 9108 4602 9188 5162
rect 9328 5202 9428 5442
rect 9328 5082 9348 5202
rect 9348 5072 9428 5082
rect 11248 5522 11348 5542
rect 11248 5422 11268 5522
rect 11328 5422 11348 5522
rect 11248 5242 11348 5422
rect 9108 4512 9188 4522
rect 10528 4822 10608 4832
rect 8808 4402 8868 4412
rect 7048 4162 7108 4172
rect 3280 2930 3400 2940
rect 4360 3100 4560 3134
rect 2920 2390 3020 2420
rect 4360 2900 4380 3100
rect 2700 2160 2760 2170
rect 2700 1990 2760 2080
rect 2920 2160 3000 2390
rect 2920 2070 3000 2080
rect 2680 1980 2760 1990
rect 2680 1910 2760 1920
rect 2040 1870 2120 1880
rect 2040 1660 2120 1670
rect 2340 1850 2480 1870
rect 2700 1860 2760 1910
rect 2460 1690 2480 1850
rect 2040 1460 2100 1660
rect 2040 1450 2140 1460
rect 2040 1250 2060 1450
rect 2040 1240 2140 1250
rect 2340 1430 2480 1690
rect 2680 1850 2760 1860
rect 2740 1670 2760 1850
rect 2680 1660 2760 1670
rect 2460 1270 2480 1430
rect 2040 1040 2100 1240
rect 2040 1030 2120 1040
rect 2040 850 2060 1030
rect 2040 840 2120 850
rect 2340 1010 2480 1270
rect 2460 850 2480 1010
rect 2040 620 2100 840
rect 2040 610 2120 620
rect 2040 430 2060 610
rect 2040 420 2120 430
rect 2340 590 2480 850
rect 2460 430 2480 590
rect 2040 350 2100 420
rect 1580 60 1700 70
rect 2340 210 2480 430
rect 2700 1450 2760 1660
rect 2700 1030 2760 1270
rect 2700 610 2760 850
rect 2700 370 2760 430
rect 2340 60 2480 70
rect 160 -1384 500 40
rect 4360 -1384 4560 2900
rect 5360 3080 5560 3100
rect 5360 2920 5380 3080
rect 5540 2920 5560 3080
rect 5360 2120 5560 2920
rect 5360 1960 5380 2120
rect 5540 1960 5560 2120
rect 7048 2102 7108 4102
rect 8388 4062 8468 4072
rect 8388 3862 8468 4002
rect 8808 4062 8868 4322
rect 9108 4282 9168 4292
rect 9168 4222 9188 4262
rect 9108 4162 9188 4222
rect 9168 4102 9188 4162
rect 9108 4082 9188 4102
rect 8808 3992 8868 4002
rect 7048 2012 7108 2022
rect 7908 3822 7988 3832
rect 5360 1940 5560 1960
rect 158 -1616 500 -1384
rect 158 -1916 198 -1616
rect 458 -1734 500 -1616
rect 4358 -1634 4560 -1384
rect 4980 1800 5140 1820
rect 4980 1640 5000 1800
rect 5120 1640 5140 1800
rect 7908 1782 7988 3742
rect 7908 1652 7988 1662
rect 8108 3802 8208 3812
rect 8448 3762 8468 3862
rect 9148 3802 9208 3812
rect 8388 3752 8448 3762
rect 8108 2682 8208 3702
rect 8848 3682 8948 3702
rect 8848 3622 8868 3682
rect 8928 3622 8948 3682
rect 8848 3122 8948 3622
rect 8848 3062 8868 3122
rect 8928 3062 8948 3122
rect 8848 3042 8948 3062
rect 9128 3622 9148 3802
rect 9208 3622 9228 3802
rect 458 -1916 498 -1734
rect 158 -1956 498 -1916
rect 4358 -2196 4558 -1634
rect 4980 -2150 5140 1640
rect 8108 -1658 8208 2602
rect 9128 2272 9228 3622
rect 10188 3562 10248 3572
rect 10248 3502 10268 3562
rect 10188 3182 10268 3502
rect 10188 3122 10208 3182
rect 9528 3102 9628 3122
rect 10208 3112 10268 3122
rect 10528 3202 10608 4742
rect 11248 4682 11268 5242
rect 11328 4682 11348 5242
rect 11248 4642 11348 4682
rect 12020 5400 12220 5420
rect 12020 5240 12040 5400
rect 12200 5240 12220 5400
rect 10588 3142 10608 3202
rect 9588 2862 9628 3102
rect 9528 2682 9628 2862
rect 9008 2262 9428 2272
rect 9008 1972 9428 1982
rect 8108 -1718 8128 -1658
rect 8188 -1718 8208 -1658
rect 8108 -1738 8208 -1718
rect 9528 -1658 9628 2602
rect 10528 2082 10608 3142
rect 12020 3240 12220 5240
rect 12020 3080 12040 3240
rect 12200 3080 12220 3240
rect 12020 3060 12220 3080
rect 10328 2062 10808 2082
rect 10328 1802 10348 2062
rect 10788 1802 10808 2062
rect 10328 1782 10808 1802
rect 12880 1780 13100 6560
rect 17320 5880 17500 5890
rect 17320 5690 17500 5700
rect 17360 5520 17460 5530
rect 17340 5440 17360 5520
rect 13080 1580 13100 1780
rect 13700 5400 13860 5420
rect 13700 5240 13720 5400
rect 13840 5240 13860 5400
rect 12880 1570 13080 1580
rect 13080 1100 13280 1120
rect 13260 920 13280 1100
rect 13080 -1384 13280 920
rect 13700 -1384 13860 5240
rect 14280 5400 14460 5420
rect 14280 5240 14300 5400
rect 14440 5240 14460 5400
rect 14280 4320 14460 5240
rect 14280 4160 14320 4320
rect 14280 4140 14460 4160
rect 15860 4380 15960 4400
rect 15940 4020 15960 4380
rect 14580 3800 14680 3810
rect 14580 3580 14680 3700
rect 15860 3800 15960 4020
rect 15940 3720 15960 3800
rect 15860 3680 15960 3720
rect 16780 3940 16860 3950
rect 14580 3180 14600 3580
rect 14660 3180 14680 3580
rect 14580 3160 14680 3180
rect 16440 3440 16560 3480
rect 16540 3220 16560 3440
rect 16440 2640 16560 3220
rect 16440 2520 16560 2540
rect 14020 1780 14160 1790
rect 14160 1580 14180 1780
rect 14020 -1384 14180 1580
rect 14300 1420 14500 1460
rect 14300 1280 14340 1420
rect 14460 1280 14500 1420
rect 14300 540 14500 1280
rect 14890 1000 14970 1010
rect 14890 920 14970 930
rect 15340 1000 15400 1010
rect 14620 840 14700 850
rect 14300 360 14340 540
rect 14460 360 14500 540
rect 14300 -1384 14500 360
rect 14600 760 14620 840
rect 14600 160 14700 760
rect 14900 730 14940 920
rect 14900 720 14960 730
rect 14900 650 14960 660
rect 15340 500 15400 940
rect 16780 960 16860 3880
rect 17180 3820 17300 3830
rect 17180 3690 17300 3700
rect 17180 2640 17260 2650
rect 17180 1860 17260 2520
rect 17240 1800 17260 1860
rect 17180 1790 17240 1800
rect 17080 1760 17140 1770
rect 16900 1710 16970 1720
rect 16900 1090 16970 1600
rect 17340 1720 17460 5440
rect 23760 2680 23980 2700
rect 23760 2500 23780 2680
rect 23960 2500 23980 2680
rect 23760 2480 23980 2500
rect 17340 1640 17360 1720
rect 17440 1640 17460 1720
rect 17340 1600 17460 1640
rect 17340 1520 17360 1600
rect 17440 1520 17460 1600
rect 17340 1460 17460 1520
rect 17340 1380 17360 1460
rect 17440 1380 17460 1460
rect 17340 1320 17460 1380
rect 17340 1240 17360 1320
rect 17440 1240 17460 1320
rect 17340 1180 17460 1240
rect 16900 1080 16980 1090
rect 16900 990 16980 1000
rect 16780 890 16860 900
rect 17080 720 17140 1180
rect 17060 710 17140 720
rect 17200 1100 17260 1110
rect 17200 780 17260 1040
rect 17200 710 17260 720
rect 17120 650 17140 710
rect 17060 640 17140 650
rect 17080 480 17140 640
rect 17320 620 17420 800
rect 15340 430 15400 440
rect 14600 10 14700 20
rect 15600 140 15940 200
rect 15600 20 15640 140
rect 15900 20 15940 140
rect 15600 -1384 15940 20
rect 17320 140 17420 480
rect 17320 10 17420 20
rect 9528 -1718 9548 -1658
rect 9608 -1718 9628 -1658
rect 9528 -1738 9628 -1718
rect 13078 -1620 13280 -1384
rect 13698 -1620 13860 -1384
rect 14018 -1620 14180 -1384
rect 14298 -1620 14500 -1384
rect 4358 -2306 4558 -2296
rect 4960 -2160 5160 -2150
rect 13078 -2176 13278 -1620
rect 13078 -2276 13098 -2176
rect 13258 -2276 13278 -2176
rect 13078 -2296 13278 -2276
rect 13698 -2196 13858 -1620
rect 13698 -2276 13718 -2196
rect 13838 -2276 13858 -2196
rect 13698 -2296 13858 -2276
rect 14018 -2176 14178 -1620
rect 14298 -2176 14498 -1620
rect 15598 -1630 15940 -1384
rect 15598 -1636 15938 -1630
rect 15598 -1876 15678 -1636
rect 15878 -1876 15938 -1636
rect 15598 -1956 15938 -1876
rect 14298 -2276 14318 -2176
rect 14478 -2276 14498 -2176
rect 14298 -2296 14498 -2276
rect 4960 -2310 5160 -2300
rect 14018 -2306 14178 -2296
<< via2 >>
rect 6940 6880 7260 7160
rect 3500 5320 4000 5480
rect 8760 5540 8960 5900
rect 9008 1982 9428 2262
rect 10348 1802 10788 2062
rect 17320 5700 17500 5880
rect 17180 3700 17300 3820
rect 23780 2500 23960 2680
rect 17320 40 17420 140
<< metal3 >>
rect 6930 7160 7270 7165
rect 6930 6880 6940 7160
rect 7260 6880 7270 7160
rect 6930 6875 7270 6880
rect 6980 5920 17520 5940
rect 6980 5720 7000 5920
rect 7260 5900 17520 5920
rect 7260 5720 8760 5900
rect 6980 5700 8760 5720
rect 8720 5540 8760 5700
rect 8960 5880 17520 5900
rect 8960 5700 17320 5880
rect 17500 5700 17520 5880
rect 8960 5540 9000 5700
rect 17310 5695 17510 5700
rect 8750 5535 8970 5540
rect 3490 5480 4010 5485
rect 3480 5320 3500 5480
rect 4000 5320 6920 5480
rect 3480 5300 6920 5320
rect 7240 5300 7250 5480
rect 3480 5280 7220 5300
rect 17160 3820 17320 3840
rect 17160 3700 17180 3820
rect 17300 3700 17320 3820
rect 17160 3680 17320 3700
rect 9008 2267 9428 2282
rect 8998 2262 9438 2267
rect 8998 1982 9008 2262
rect 9428 1982 9438 2262
rect 8998 1977 9438 1982
rect 10328 2062 10808 2082
rect 9008 1502 9428 1977
rect 10328 1802 10348 2062
rect 10788 1802 10808 2062
rect 10328 1782 10808 1802
rect 5368 1474 11740 1502
rect 5368 -1550 11656 1474
rect 11720 -1550 11740 1474
rect 17720 160 23240 5852
rect 23760 2680 23980 2700
rect 23760 2500 23780 2680
rect 23960 2500 23980 2680
rect 23760 2480 23980 2500
rect 24100 160 29620 5852
rect 17280 140 29620 160
rect 17280 40 17320 140
rect 17420 124 29620 140
rect 17420 60 17748 124
rect 23212 60 24128 124
rect 29592 60 29620 124
rect 17420 40 29620 60
rect 17280 0 24580 40
rect 5368 -1578 11740 -1550
<< via3 >>
rect 6940 6880 7260 7160
rect 7000 5720 7260 5920
rect 6920 5300 7240 5480
rect 17180 3700 17300 3820
rect 10348 1802 10788 2062
rect 11656 -1550 11720 1474
rect 23780 2500 23960 2680
rect 17748 60 23212 124
rect 24128 60 29592 124
<< mimcap >>
rect 17760 5772 23200 5812
rect 5408 1422 11408 1462
rect 5408 -1498 5448 1422
rect 11368 -1498 11408 1422
rect 17760 412 17800 5772
rect 23160 412 23200 5772
rect 17760 372 23200 412
rect 24140 5772 29580 5812
rect 24140 412 24180 5772
rect 29540 412 29580 5772
rect 24140 372 29580 412
rect 5408 -1538 11408 -1498
<< mimcapcontact >>
rect 5448 -1498 11368 1422
rect 17800 412 23160 5772
rect 24180 412 29540 5772
<< metal4 >>
rect 6900 7160 7280 7240
rect 6900 6880 6940 7160
rect 7260 6880 7280 7160
rect 6900 6401 7280 6880
rect 6899 6279 7280 6401
rect 6900 5920 7280 6279
rect 6900 5720 7000 5920
rect 7260 5720 7280 5920
rect 6900 5480 7280 5720
rect 6900 5300 6920 5480
rect 7240 5300 7280 5480
rect 6900 5150 7280 5300
rect 17799 5772 23161 5773
rect 17799 3840 17800 5772
rect 16940 3820 17800 3840
rect 16940 3700 17180 3820
rect 17300 3700 17800 3820
rect 16940 3400 17800 3700
rect 10328 2062 10808 2082
rect 10328 1802 10348 2062
rect 10788 1802 10808 2062
rect 10328 1782 10808 1802
rect 10348 1423 10788 1782
rect 11640 1474 11736 1490
rect 5447 1422 11369 1423
rect 5447 -1498 5448 1422
rect 11368 -1498 11369 1422
rect 5447 -1499 11369 -1498
rect 11640 -1550 11656 1474
rect 11720 -1550 11736 1474
rect 17799 412 17800 3400
rect 23160 412 23161 5772
rect 24179 5772 29541 5773
rect 24179 2800 24180 5772
rect 23920 2700 24180 2800
rect 23760 2680 24180 2700
rect 23760 2500 23780 2680
rect 23960 2500 24180 2680
rect 23760 2480 24180 2500
rect 23920 2360 24180 2480
rect 17799 411 23161 412
rect 24179 412 24180 2360
rect 29540 412 29541 5772
rect 24179 411 29541 412
rect 17732 124 23228 140
rect 17732 60 17748 124
rect 23212 60 23228 124
rect 17732 44 23228 60
rect 24112 124 29608 140
rect 24112 60 24128 124
rect 29592 60 29608 124
rect 24112 44 29608 60
rect 11640 -1566 11736 -1550
<< comment >>
rect 17700 20 17720 40
rect 24080 20 24100 40
rect 23600 0 23620 20
rect -20 -20 0 0
rect 14280 -20 14300 0
rect 5340 -1820 5360 -1800
<< labels >>
flabel metal1 4306 3508 4334 3538 0 FreeSans 1600 0 0 0 vtd
flabel metal1 11842 6654 11886 6698 0 FreeSans 800 0 0 0 out_sigma
flabel metal1 -62 -1956 138 -1756 0 FreeSans 1600 0 0 0 gnd
port 1 nsew
flabel metal1 14278 -2576 14478 -2376 0 FreeSans 1600 0 0 0 vpwr
port 4 nsew
flabel metal1 13078 -2576 13278 -2376 0 FreeSans 1600 0 0 0 clk
port 2 nsew
flabel metal1 13658 -2576 13858 -2376 0 FreeSans 1600 0 0 0 out_buff
port 7 nsew
flabel metal1 14018 -2576 14218 -2376 0 FreeSans 1600 0 0 0 out_sigma
port 9 nsew
flabel metal1 4958 -2576 5158 -2376 0 FreeSans 1600 0 0 0 ib
port 5 nsew
flabel metal1 4360 -2580 4560 -2380 0 FreeSans 1600 0 0 0 vts
port 8 nsew
flabel metal1 200 6580 400 6780 0 FreeSans 1600 0 0 0 out
port 3 nsew
flabel metal1 6980 7340 7180 7540 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 14300 1260 14500 1460 0 FreeSans 1600 0 0 0 sigma-delta_0.vpwr
flabel metal1 14300 920 14500 1120 0 FreeSans 1600 0 0 0 sigma-delta_0.clk
flabel metal1 14300 360 14500 560 0 FreeSans 1600 0 0 0 sigma-delta_0.reset_b_dff
flabel metal1 15720 0 15920 200 0 FreeSans 1600 0 0 0 sigma-delta_0.gnd
flabel metal1 17340 5680 17540 5880 0 FreeSans 1600 0 0 0 sigma-delta_0.vd
flabel metal1 16080 3740 16140 3760 0 FreeSans 800 0 0 0 sigma-delta_0.in_int
flabel metal1 16140 3340 16200 3360 0 FreeSans 800 0 0 0 sigma-delta_0.in_comp
flabel metal1 14300 1560 14500 1760 0 FreeSans 1600 0 0 0 sigma-delta_0.out
flabel metal1 14300 4140 14500 4340 0 FreeSans 1600 0 0 0 sigma-delta_0.in
flabel locali 16352 1026 16381 1061 0 FreeSans 200 0 0 0 sigma-delta_0.x1.Q
flabel locali 16654 1029 16676 1062 0 FreeSans 200 0 0 0 sigma-delta_0.x1.Q_N
flabel locali 16079 961 16113 995 0 FreeSans 400 0 0 0 sigma-delta_0.x1.RESET_B
flabel locali 14903 1097 14937 1131 0 FreeSans 400 0 0 0 sigma-delta_0.x1.D
flabel locali 14628 1097 14662 1131 0 FreeSans 400 0 0 0 sigma-delta_0.x1.CLK
flabel locali 14628 1029 14662 1063 0 FreeSans 400 0 0 0 sigma-delta_0.x1.CLK
flabel locali 16079 1029 16113 1063 0 FreeSans 400 0 0 0 sigma-delta_0.x1.RESET_B
flabel metal1 14627 791 14661 825 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VGND
flabel metal1 14627 1335 14661 1369 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VPWR
flabel nwell 14627 1335 14661 1369 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VPB
flabel pwell 14627 791 14661 825 0 FreeSans 200 0 0 0 sigma-delta_0.x1.VNB
rlabel comment 14598 808 14598 808 4 sigma-delta_0.x1.dfrbp_1
rlabel locali 16079 935 16127 1015 1 sigma-delta_0.x1.RESET_B
rlabel locali 16019 1015 16127 1089 1 sigma-delta_0.x1.RESET_B
rlabel metal1 16067 955 16125 964 1 sigma-delta_0.x1.RESET_B
rlabel metal1 16007 1001 16065 1064 1 sigma-delta_0.x1.RESET_B
rlabel metal1 16007 992 16125 1001 1 sigma-delta_0.x1.RESET_B
rlabel metal1 15347 992 15477 1001 1 sigma-delta_0.x1.RESET_B
rlabel metal1 15347 964 16125 992 1 sigma-delta_0.x1.RESET_B
rlabel metal1 15347 955 15477 964 1 sigma-delta_0.x1.RESET_B
rlabel metal1 14598 760 16714 856 1 sigma-delta_0.x1.VGND
rlabel metal1 14598 1304 16714 1400 1 sigma-delta_0.x1.VPWR
flabel metal1 480 5300 680 5500 0 FreeSans 256 0 0 0 sensor_0.vd
flabel metal1 160 0 360 200 0 FreeSans 256 0 0 0 sensor_0.gnd
flabel metal1 4040 2900 4240 3100 0 FreeSans 256 0 0 0 sensor_0.vts
flabel metal1 4040 3360 4240 3560 0 FreeSans 256 0 0 0 sensor_0.vtd
flabel metal2 860 3580 880 3600 0 FreeSans 800 0 0 0 sensor_0.a
flabel metal2 2380 4440 2400 4460 0 FreeSans 800 0 0 0 sensor_0.d
flabel metal1 2500 3940 2520 3980 0 FreeSans 800 0 0 0 sensor_0.c
flabel metal2 2960 2220 2960 2240 0 FreeSans 800 0 0 0 sensor_0.b
flabel metal2 8488 4842 8508 4882 0 FreeSans 800 0 0 0 buffer_0.a
flabel metal2 9128 4842 9168 4862 0 FreeSans 800 0 0 0 buffer_0.b
flabel metal1 8748 5542 8948 5742 0 FreeSans 256 0 0 0 buffer_0.vd
flabel metal1 8568 4022 8588 4042 0 FreeSans 800 0 0 0 buffer_0.c
flabel metal1 5368 1622 5568 1822 0 FreeSans 256 0 0 0 buffer_0.ib
flabel metal1 5368 1942 5568 2142 0 FreeSans 256 0 0 0 buffer_0.in
flabel metal1 7188 3102 7208 3122 0 FreeSans 800 0 0 0 buffer_0.d
flabel metal1 12028 3062 12228 3262 0 FreeSans 256 0 0 0 buffer_0.out
flabel metal1 5368 -1798 5568 -1598 0 FreeSans 256 0 0 0 buffer_0.gnd
<< end >>
