magic
tech sky130A
magscale 1 2
timestamp 1645148224
<< metal4 >>
rect -2329 6809 2329 6850
rect -2329 2391 2073 6809
rect 2309 2391 2329 6809
rect -2329 2350 2329 2391
rect -2329 2209 2329 2250
rect -2329 -2209 2073 2209
rect 2309 -2209 2329 2209
rect -2329 -2250 2329 -2209
rect -2329 -2391 2329 -2350
rect -2329 -6809 2073 -2391
rect 2309 -6809 2329 -2391
rect -2329 -6850 2329 -6809
<< via4 >>
rect 2073 2391 2309 6809
rect 2073 -2209 2309 2209
rect 2073 -6809 2309 -2391
<< mimcap2 >>
rect -2229 6710 2071 6750
rect -2229 2490 -1767 6710
rect 1609 2490 2071 6710
rect -2229 2450 2071 2490
rect -2229 2110 2071 2150
rect -2229 -2110 -1767 2110
rect 1609 -2110 2071 2110
rect -2229 -2150 2071 -2110
rect -2229 -2490 2071 -2450
rect -2229 -6710 -1767 -2490
rect 1609 -6710 2071 -2490
rect -2229 -6750 2071 -6710
<< mimcap2contact >>
rect -1767 2490 1609 6710
rect -1767 -2110 1609 2110
rect -1767 -6710 1609 -2490
<< metal5 >>
rect -239 6734 81 6900
rect 2031 6809 2351 6900
rect -1791 6710 1633 6734
rect -1791 2490 -1767 6710
rect 1609 2490 1633 6710
rect -1791 2466 1633 2490
rect -239 2134 81 2466
rect 2031 2391 2073 6809
rect 2309 2391 2351 6809
rect 2031 2209 2351 2391
rect -1791 2110 1633 2134
rect -1791 -2110 -1767 2110
rect 1609 -2110 1633 2110
rect -1791 -2134 1633 -2110
rect -239 -2466 81 -2134
rect 2031 -2209 2073 2209
rect 2309 -2209 2351 2209
rect 2031 -2391 2351 -2209
rect -1791 -2490 1633 -2466
rect -1791 -6710 -1767 -2490
rect 1609 -6710 1633 -2490
rect -1791 -6734 1633 -6710
rect -239 -6900 81 -6734
rect 2031 -6809 2073 -2391
rect 2309 -6809 2351 -2391
rect 2031 -6900 2351 -6809
<< properties >>
string FIXED_BBOX -2329 2350 2171 6850
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 21.5 l 21.5 val 940.84 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
