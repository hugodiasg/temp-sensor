magic
tech sky130A
timestamp 1645729143
<< metal4 >>
rect 19400 21490 21500 21500
rect 19400 20910 20910 21490
rect 21490 20910 21500 21490
rect 19400 20900 21500 20910
<< via4 >>
rect 20910 20910 21490 21490
<< metal5 >>
rect 20000 34400 35000 35000
rect 20000 33500 34100 34100
rect 20000 20600 20600 33500
rect 20898 21500 21502 21502
rect 33500 21500 34100 33500
rect 20898 21490 34100 21500
rect 20898 20910 20910 21490
rect 21490 20910 34100 21490
rect 20898 20900 34100 20910
rect 20898 20898 21502 20900
rect 34400 20600 35000 34400
rect 20000 20000 35000 20600
<< end >>
