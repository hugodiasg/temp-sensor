magic
tech sky130A
timestamp 1643668240
<< metal3 >>
rect 7000 -500 7500 6900
<< metal4 >>
rect 0 13400 13900 13900
rect 0 12600 13100 13100
rect 0 500 500 12600
rect 800 11800 12300 12300
rect 800 1300 1300 11800
rect 1600 11000 11500 11500
rect 1600 2100 2100 11000
rect 2400 10200 10700 10700
rect 2400 2900 2900 10200
rect 3200 9400 9900 9900
rect 3200 3700 3700 9400
rect 4000 8600 9100 9100
rect 4000 4500 4500 8600
rect 4800 7800 8300 8300
rect 4800 5300 5300 7800
rect 5600 7000 7500 7500
rect 5600 6100 6100 7000
rect 7000 6400 7500 7000
rect 7800 6100 8300 7800
rect 5600 5600 8300 6100
rect 8600 5300 9100 8600
rect 4800 4800 9100 5300
rect 9400 4500 9900 9400
rect 4000 4000 9900 4500
rect 10200 3700 10700 10200
rect 3200 3200 10700 3700
rect 11000 2900 11500 11000
rect 2400 2400 11500 2900
rect 11800 2100 12300 11800
rect 1600 1600 12300 2100
rect 12600 1300 13100 12600
rect 800 800 13100 1300
rect 13400 500 13900 13400
rect 0 0 13900 500
<< end >>
