magic
tech sky130A
timestamp 1700063261
<< nmos >>
rect -1340 -50 -1240 50
rect -1211 -50 -1111 50
rect -1082 -50 -982 50
rect -953 -50 -853 50
rect -824 -50 -724 50
rect -695 -50 -595 50
rect -566 -50 -466 50
rect -437 -50 -337 50
rect -308 -50 -208 50
rect -179 -50 -79 50
rect -50 -50 50 50
rect 79 -50 179 50
rect 208 -50 308 50
rect 337 -50 437 50
rect 466 -50 566 50
rect 595 -50 695 50
rect 724 -50 824 50
rect 853 -50 953 50
rect 982 -50 1082 50
rect 1111 -50 1211 50
rect 1240 -50 1340 50
<< ndiff >>
rect -1369 44 -1340 50
rect -1369 -44 -1363 44
rect -1346 -44 -1340 44
rect -1369 -50 -1340 -44
rect -1240 44 -1211 50
rect -1240 -44 -1234 44
rect -1217 -44 -1211 44
rect -1240 -50 -1211 -44
rect -1111 44 -1082 50
rect -1111 -44 -1105 44
rect -1088 -44 -1082 44
rect -1111 -50 -1082 -44
rect -982 44 -953 50
rect -982 -44 -976 44
rect -959 -44 -953 44
rect -982 -50 -953 -44
rect -853 44 -824 50
rect -853 -44 -847 44
rect -830 -44 -824 44
rect -853 -50 -824 -44
rect -724 44 -695 50
rect -724 -44 -718 44
rect -701 -44 -695 44
rect -724 -50 -695 -44
rect -595 44 -566 50
rect -595 -44 -589 44
rect -572 -44 -566 44
rect -595 -50 -566 -44
rect -466 44 -437 50
rect -466 -44 -460 44
rect -443 -44 -437 44
rect -466 -50 -437 -44
rect -337 44 -308 50
rect -337 -44 -331 44
rect -314 -44 -308 44
rect -337 -50 -308 -44
rect -208 44 -179 50
rect -208 -44 -202 44
rect -185 -44 -179 44
rect -208 -50 -179 -44
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
rect 179 44 208 50
rect 179 -44 185 44
rect 202 -44 208 44
rect 179 -50 208 -44
rect 308 44 337 50
rect 308 -44 314 44
rect 331 -44 337 44
rect 308 -50 337 -44
rect 437 44 466 50
rect 437 -44 443 44
rect 460 -44 466 44
rect 437 -50 466 -44
rect 566 44 595 50
rect 566 -44 572 44
rect 589 -44 595 44
rect 566 -50 595 -44
rect 695 44 724 50
rect 695 -44 701 44
rect 718 -44 724 44
rect 695 -50 724 -44
rect 824 44 853 50
rect 824 -44 830 44
rect 847 -44 853 44
rect 824 -50 853 -44
rect 953 44 982 50
rect 953 -44 959 44
rect 976 -44 982 44
rect 953 -50 982 -44
rect 1082 44 1111 50
rect 1082 -44 1088 44
rect 1105 -44 1111 44
rect 1082 -50 1111 -44
rect 1211 44 1240 50
rect 1211 -44 1217 44
rect 1234 -44 1240 44
rect 1211 -50 1240 -44
rect 1340 44 1369 50
rect 1340 -44 1346 44
rect 1363 -44 1369 44
rect 1340 -50 1369 -44
<< ndiffc >>
rect -1363 -44 -1346 44
rect -1234 -44 -1217 44
rect -1105 -44 -1088 44
rect -976 -44 -959 44
rect -847 -44 -830 44
rect -718 -44 -701 44
rect -589 -44 -572 44
rect -460 -44 -443 44
rect -331 -44 -314 44
rect -202 -44 -185 44
rect -73 -44 -56 44
rect 56 -44 73 44
rect 185 -44 202 44
rect 314 -44 331 44
rect 443 -44 460 44
rect 572 -44 589 44
rect 701 -44 718 44
rect 830 -44 847 44
rect 959 -44 976 44
rect 1088 -44 1105 44
rect 1217 -44 1234 44
rect 1346 -44 1363 44
<< poly >>
rect -1340 86 -1240 94
rect -1340 69 -1332 86
rect -1248 69 -1240 86
rect -1340 50 -1240 69
rect -1211 86 -1111 94
rect -1211 69 -1203 86
rect -1119 69 -1111 86
rect -1211 50 -1111 69
rect -1082 86 -982 94
rect -1082 69 -1074 86
rect -990 69 -982 86
rect -1082 50 -982 69
rect -953 86 -853 94
rect -953 69 -945 86
rect -861 69 -853 86
rect -953 50 -853 69
rect -824 86 -724 94
rect -824 69 -816 86
rect -732 69 -724 86
rect -824 50 -724 69
rect -695 86 -595 94
rect -695 69 -687 86
rect -603 69 -595 86
rect -695 50 -595 69
rect -566 86 -466 94
rect -566 69 -558 86
rect -474 69 -466 86
rect -566 50 -466 69
rect -437 86 -337 94
rect -437 69 -429 86
rect -345 69 -337 86
rect -437 50 -337 69
rect -308 86 -208 94
rect -308 69 -300 86
rect -216 69 -208 86
rect -308 50 -208 69
rect -179 86 -79 94
rect -179 69 -171 86
rect -87 69 -79 86
rect -179 50 -79 69
rect -50 86 50 94
rect -50 69 -42 86
rect 42 69 50 86
rect -50 50 50 69
rect 79 86 179 94
rect 79 69 87 86
rect 171 69 179 86
rect 79 50 179 69
rect 208 86 308 94
rect 208 69 216 86
rect 300 69 308 86
rect 208 50 308 69
rect 337 86 437 94
rect 337 69 345 86
rect 429 69 437 86
rect 337 50 437 69
rect 466 86 566 94
rect 466 69 474 86
rect 558 69 566 86
rect 466 50 566 69
rect 595 86 695 94
rect 595 69 603 86
rect 687 69 695 86
rect 595 50 695 69
rect 724 86 824 94
rect 724 69 732 86
rect 816 69 824 86
rect 724 50 824 69
rect 853 86 953 94
rect 853 69 861 86
rect 945 69 953 86
rect 853 50 953 69
rect 982 86 1082 94
rect 982 69 990 86
rect 1074 69 1082 86
rect 982 50 1082 69
rect 1111 86 1211 94
rect 1111 69 1119 86
rect 1203 69 1211 86
rect 1111 50 1211 69
rect 1240 86 1340 94
rect 1240 69 1248 86
rect 1332 69 1340 86
rect 1240 50 1340 69
rect -1340 -69 -1240 -50
rect -1340 -86 -1332 -69
rect -1248 -86 -1240 -69
rect -1340 -94 -1240 -86
rect -1211 -69 -1111 -50
rect -1211 -86 -1203 -69
rect -1119 -86 -1111 -69
rect -1211 -94 -1111 -86
rect -1082 -69 -982 -50
rect -1082 -86 -1074 -69
rect -990 -86 -982 -69
rect -1082 -94 -982 -86
rect -953 -69 -853 -50
rect -953 -86 -945 -69
rect -861 -86 -853 -69
rect -953 -94 -853 -86
rect -824 -69 -724 -50
rect -824 -86 -816 -69
rect -732 -86 -724 -69
rect -824 -94 -724 -86
rect -695 -69 -595 -50
rect -695 -86 -687 -69
rect -603 -86 -595 -69
rect -695 -94 -595 -86
rect -566 -69 -466 -50
rect -566 -86 -558 -69
rect -474 -86 -466 -69
rect -566 -94 -466 -86
rect -437 -69 -337 -50
rect -437 -86 -429 -69
rect -345 -86 -337 -69
rect -437 -94 -337 -86
rect -308 -69 -208 -50
rect -308 -86 -300 -69
rect -216 -86 -208 -69
rect -308 -94 -208 -86
rect -179 -69 -79 -50
rect -179 -86 -171 -69
rect -87 -86 -79 -69
rect -179 -94 -79 -86
rect -50 -69 50 -50
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -50 -94 50 -86
rect 79 -69 179 -50
rect 79 -86 87 -69
rect 171 -86 179 -69
rect 79 -94 179 -86
rect 208 -69 308 -50
rect 208 -86 216 -69
rect 300 -86 308 -69
rect 208 -94 308 -86
rect 337 -69 437 -50
rect 337 -86 345 -69
rect 429 -86 437 -69
rect 337 -94 437 -86
rect 466 -69 566 -50
rect 466 -86 474 -69
rect 558 -86 566 -69
rect 466 -94 566 -86
rect 595 -69 695 -50
rect 595 -86 603 -69
rect 687 -86 695 -69
rect 595 -94 695 -86
rect 724 -69 824 -50
rect 724 -86 732 -69
rect 816 -86 824 -69
rect 724 -94 824 -86
rect 853 -69 953 -50
rect 853 -86 861 -69
rect 945 -86 953 -69
rect 853 -94 953 -86
rect 982 -69 1082 -50
rect 982 -86 990 -69
rect 1074 -86 1082 -69
rect 982 -94 1082 -86
rect 1111 -69 1211 -50
rect 1111 -86 1119 -69
rect 1203 -86 1211 -69
rect 1111 -94 1211 -86
rect 1240 -69 1340 -50
rect 1240 -86 1248 -69
rect 1332 -86 1340 -69
rect 1240 -94 1340 -86
<< polycont >>
rect -1332 69 -1248 86
rect -1203 69 -1119 86
rect -1074 69 -990 86
rect -945 69 -861 86
rect -816 69 -732 86
rect -687 69 -603 86
rect -558 69 -474 86
rect -429 69 -345 86
rect -300 69 -216 86
rect -171 69 -87 86
rect -42 69 42 86
rect 87 69 171 86
rect 216 69 300 86
rect 345 69 429 86
rect 474 69 558 86
rect 603 69 687 86
rect 732 69 816 86
rect 861 69 945 86
rect 990 69 1074 86
rect 1119 69 1203 86
rect 1248 69 1332 86
rect -1332 -86 -1248 -69
rect -1203 -86 -1119 -69
rect -1074 -86 -990 -69
rect -945 -86 -861 -69
rect -816 -86 -732 -69
rect -687 -86 -603 -69
rect -558 -86 -474 -69
rect -429 -86 -345 -69
rect -300 -86 -216 -69
rect -171 -86 -87 -69
rect -42 -86 42 -69
rect 87 -86 171 -69
rect 216 -86 300 -69
rect 345 -86 429 -69
rect 474 -86 558 -69
rect 603 -86 687 -69
rect 732 -86 816 -69
rect 861 -86 945 -69
rect 990 -86 1074 -69
rect 1119 -86 1203 -69
rect 1248 -86 1332 -69
<< locali >>
rect -1340 69 -1332 86
rect -1248 69 -1240 86
rect -1211 69 -1203 86
rect -1119 69 -1111 86
rect -1082 69 -1074 86
rect -990 69 -982 86
rect -953 69 -945 86
rect -861 69 -853 86
rect -824 69 -816 86
rect -732 69 -724 86
rect -695 69 -687 86
rect -603 69 -595 86
rect -566 69 -558 86
rect -474 69 -466 86
rect -437 69 -429 86
rect -345 69 -337 86
rect -308 69 -300 86
rect -216 69 -208 86
rect -179 69 -171 86
rect -87 69 -79 86
rect -50 69 -42 86
rect 42 69 50 86
rect 79 69 87 86
rect 171 69 179 86
rect 208 69 216 86
rect 300 69 308 86
rect 337 69 345 86
rect 429 69 437 86
rect 466 69 474 86
rect 558 69 566 86
rect 595 69 603 86
rect 687 69 695 86
rect 724 69 732 86
rect 816 69 824 86
rect 853 69 861 86
rect 945 69 953 86
rect 982 69 990 86
rect 1074 69 1082 86
rect 1111 69 1119 86
rect 1203 69 1211 86
rect 1240 69 1248 86
rect 1332 69 1340 86
rect -1363 44 -1346 52
rect -1363 -52 -1346 -44
rect -1234 44 -1217 52
rect -1234 -52 -1217 -44
rect -1105 44 -1088 52
rect -1105 -52 -1088 -44
rect -976 44 -959 52
rect -976 -52 -959 -44
rect -847 44 -830 52
rect -847 -52 -830 -44
rect -718 44 -701 52
rect -718 -52 -701 -44
rect -589 44 -572 52
rect -589 -52 -572 -44
rect -460 44 -443 52
rect -460 -52 -443 -44
rect -331 44 -314 52
rect -331 -52 -314 -44
rect -202 44 -185 52
rect -202 -52 -185 -44
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect 185 44 202 52
rect 185 -52 202 -44
rect 314 44 331 52
rect 314 -52 331 -44
rect 443 44 460 52
rect 443 -52 460 -44
rect 572 44 589 52
rect 572 -52 589 -44
rect 701 44 718 52
rect 701 -52 718 -44
rect 830 44 847 52
rect 830 -52 847 -44
rect 959 44 976 52
rect 959 -52 976 -44
rect 1088 44 1105 52
rect 1088 -52 1105 -44
rect 1217 44 1234 52
rect 1217 -52 1234 -44
rect 1346 44 1363 52
rect 1346 -52 1363 -44
rect -1340 -86 -1332 -69
rect -1248 -86 -1240 -69
rect -1211 -86 -1203 -69
rect -1119 -86 -1111 -69
rect -1082 -86 -1074 -69
rect -990 -86 -982 -69
rect -953 -86 -945 -69
rect -861 -86 -853 -69
rect -824 -86 -816 -69
rect -732 -86 -724 -69
rect -695 -86 -687 -69
rect -603 -86 -595 -69
rect -566 -86 -558 -69
rect -474 -86 -466 -69
rect -437 -86 -429 -69
rect -345 -86 -337 -69
rect -308 -86 -300 -69
rect -216 -86 -208 -69
rect -179 -86 -171 -69
rect -87 -86 -79 -69
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect 79 -86 87 -69
rect 171 -86 179 -69
rect 208 -86 216 -69
rect 300 -86 308 -69
rect 337 -86 345 -69
rect 429 -86 437 -69
rect 466 -86 474 -69
rect 558 -86 566 -69
rect 595 -86 603 -69
rect 687 -86 695 -69
rect 724 -86 732 -69
rect 816 -86 824 -69
rect 853 -86 861 -69
rect 945 -86 953 -69
rect 982 -86 990 -69
rect 1074 -86 1082 -69
rect 1111 -86 1119 -69
rect 1203 -86 1211 -69
rect 1240 -86 1248 -69
rect 1332 -86 1340 -69
<< viali >>
rect -1332 69 -1248 86
rect -1203 69 -1119 86
rect -1074 69 -990 86
rect -945 69 -861 86
rect -816 69 -732 86
rect -687 69 -603 86
rect -558 69 -474 86
rect -429 69 -345 86
rect -300 69 -216 86
rect -171 69 -87 86
rect -42 69 42 86
rect 87 69 171 86
rect 216 69 300 86
rect 345 69 429 86
rect 474 69 558 86
rect 603 69 687 86
rect 732 69 816 86
rect 861 69 945 86
rect 990 69 1074 86
rect 1119 69 1203 86
rect 1248 69 1332 86
rect -1363 -44 -1346 44
rect -1234 -44 -1217 44
rect -1105 -44 -1088 44
rect -976 -44 -959 44
rect -847 -44 -830 44
rect -718 -44 -701 44
rect -589 -44 -572 44
rect -460 -44 -443 44
rect -331 -44 -314 44
rect -202 -44 -185 44
rect -73 -44 -56 44
rect 56 -44 73 44
rect 185 -44 202 44
rect 314 -44 331 44
rect 443 -44 460 44
rect 572 -44 589 44
rect 701 -44 718 44
rect 830 -44 847 44
rect 959 -44 976 44
rect 1088 -44 1105 44
rect 1217 -44 1234 44
rect 1346 -44 1363 44
rect -1332 -86 -1248 -69
rect -1203 -86 -1119 -69
rect -1074 -86 -990 -69
rect -945 -86 -861 -69
rect -816 -86 -732 -69
rect -687 -86 -603 -69
rect -558 -86 -474 -69
rect -429 -86 -345 -69
rect -300 -86 -216 -69
rect -171 -86 -87 -69
rect -42 -86 42 -69
rect 87 -86 171 -69
rect 216 -86 300 -69
rect 345 -86 429 -69
rect 474 -86 558 -69
rect 603 -86 687 -69
rect 732 -86 816 -69
rect 861 -86 945 -69
rect 990 -86 1074 -69
rect 1119 -86 1203 -69
rect 1248 -86 1332 -69
<< metal1 >>
rect -1338 86 -1242 89
rect -1338 69 -1332 86
rect -1248 69 -1242 86
rect -1338 66 -1242 69
rect -1209 86 -1113 89
rect -1209 69 -1203 86
rect -1119 69 -1113 86
rect -1209 66 -1113 69
rect -1080 86 -984 89
rect -1080 69 -1074 86
rect -990 69 -984 86
rect -1080 66 -984 69
rect -951 86 -855 89
rect -951 69 -945 86
rect -861 69 -855 86
rect -951 66 -855 69
rect -822 86 -726 89
rect -822 69 -816 86
rect -732 69 -726 86
rect -822 66 -726 69
rect -693 86 -597 89
rect -693 69 -687 86
rect -603 69 -597 86
rect -693 66 -597 69
rect -564 86 -468 89
rect -564 69 -558 86
rect -474 69 -468 86
rect -564 66 -468 69
rect -435 86 -339 89
rect -435 69 -429 86
rect -345 69 -339 86
rect -435 66 -339 69
rect -306 86 -210 89
rect -306 69 -300 86
rect -216 69 -210 86
rect -306 66 -210 69
rect -177 86 -81 89
rect -177 69 -171 86
rect -87 69 -81 86
rect -177 66 -81 69
rect -48 86 48 89
rect -48 69 -42 86
rect 42 69 48 86
rect -48 66 48 69
rect 81 86 177 89
rect 81 69 87 86
rect 171 69 177 86
rect 81 66 177 69
rect 210 86 306 89
rect 210 69 216 86
rect 300 69 306 86
rect 210 66 306 69
rect 339 86 435 89
rect 339 69 345 86
rect 429 69 435 86
rect 339 66 435 69
rect 468 86 564 89
rect 468 69 474 86
rect 558 69 564 86
rect 468 66 564 69
rect 597 86 693 89
rect 597 69 603 86
rect 687 69 693 86
rect 597 66 693 69
rect 726 86 822 89
rect 726 69 732 86
rect 816 69 822 86
rect 726 66 822 69
rect 855 86 951 89
rect 855 69 861 86
rect 945 69 951 86
rect 855 66 951 69
rect 984 86 1080 89
rect 984 69 990 86
rect 1074 69 1080 86
rect 984 66 1080 69
rect 1113 86 1209 89
rect 1113 69 1119 86
rect 1203 69 1209 86
rect 1113 66 1209 69
rect 1242 86 1338 89
rect 1242 69 1248 86
rect 1332 69 1338 86
rect 1242 66 1338 69
rect -1366 44 -1343 50
rect -1366 -44 -1363 44
rect -1346 -44 -1343 44
rect -1366 -50 -1343 -44
rect -1237 44 -1214 50
rect -1237 -44 -1234 44
rect -1217 -44 -1214 44
rect -1237 -50 -1214 -44
rect -1108 44 -1085 50
rect -1108 -44 -1105 44
rect -1088 -44 -1085 44
rect -1108 -50 -1085 -44
rect -979 44 -956 50
rect -979 -44 -976 44
rect -959 -44 -956 44
rect -979 -50 -956 -44
rect -850 44 -827 50
rect -850 -44 -847 44
rect -830 -44 -827 44
rect -850 -50 -827 -44
rect -721 44 -698 50
rect -721 -44 -718 44
rect -701 -44 -698 44
rect -721 -50 -698 -44
rect -592 44 -569 50
rect -592 -44 -589 44
rect -572 -44 -569 44
rect -592 -50 -569 -44
rect -463 44 -440 50
rect -463 -44 -460 44
rect -443 -44 -440 44
rect -463 -50 -440 -44
rect -334 44 -311 50
rect -334 -44 -331 44
rect -314 -44 -311 44
rect -334 -50 -311 -44
rect -205 44 -182 50
rect -205 -44 -202 44
rect -185 -44 -182 44
rect -205 -50 -182 -44
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect 182 44 205 50
rect 182 -44 185 44
rect 202 -44 205 44
rect 182 -50 205 -44
rect 311 44 334 50
rect 311 -44 314 44
rect 331 -44 334 44
rect 311 -50 334 -44
rect 440 44 463 50
rect 440 -44 443 44
rect 460 -44 463 44
rect 440 -50 463 -44
rect 569 44 592 50
rect 569 -44 572 44
rect 589 -44 592 44
rect 569 -50 592 -44
rect 698 44 721 50
rect 698 -44 701 44
rect 718 -44 721 44
rect 698 -50 721 -44
rect 827 44 850 50
rect 827 -44 830 44
rect 847 -44 850 44
rect 827 -50 850 -44
rect 956 44 979 50
rect 956 -44 959 44
rect 976 -44 979 44
rect 956 -50 979 -44
rect 1085 44 1108 50
rect 1085 -44 1088 44
rect 1105 -44 1108 44
rect 1085 -50 1108 -44
rect 1214 44 1237 50
rect 1214 -44 1217 44
rect 1234 -44 1237 44
rect 1214 -50 1237 -44
rect 1343 44 1366 50
rect 1343 -44 1346 44
rect 1363 -44 1366 44
rect 1343 -50 1366 -44
rect -1338 -69 -1242 -66
rect -1338 -86 -1332 -69
rect -1248 -86 -1242 -69
rect -1338 -89 -1242 -86
rect -1209 -69 -1113 -66
rect -1209 -86 -1203 -69
rect -1119 -86 -1113 -69
rect -1209 -89 -1113 -86
rect -1080 -69 -984 -66
rect -1080 -86 -1074 -69
rect -990 -86 -984 -69
rect -1080 -89 -984 -86
rect -951 -69 -855 -66
rect -951 -86 -945 -69
rect -861 -86 -855 -69
rect -951 -89 -855 -86
rect -822 -69 -726 -66
rect -822 -86 -816 -69
rect -732 -86 -726 -69
rect -822 -89 -726 -86
rect -693 -69 -597 -66
rect -693 -86 -687 -69
rect -603 -86 -597 -69
rect -693 -89 -597 -86
rect -564 -69 -468 -66
rect -564 -86 -558 -69
rect -474 -86 -468 -69
rect -564 -89 -468 -86
rect -435 -69 -339 -66
rect -435 -86 -429 -69
rect -345 -86 -339 -69
rect -435 -89 -339 -86
rect -306 -69 -210 -66
rect -306 -86 -300 -69
rect -216 -86 -210 -69
rect -306 -89 -210 -86
rect -177 -69 -81 -66
rect -177 -86 -171 -69
rect -87 -86 -81 -69
rect -177 -89 -81 -86
rect -48 -69 48 -66
rect -48 -86 -42 -69
rect 42 -86 48 -69
rect -48 -89 48 -86
rect 81 -69 177 -66
rect 81 -86 87 -69
rect 171 -86 177 -69
rect 81 -89 177 -86
rect 210 -69 306 -66
rect 210 -86 216 -69
rect 300 -86 306 -69
rect 210 -89 306 -86
rect 339 -69 435 -66
rect 339 -86 345 -69
rect 429 -86 435 -69
rect 339 -89 435 -86
rect 468 -69 564 -66
rect 468 -86 474 -69
rect 558 -86 564 -69
rect 468 -89 564 -86
rect 597 -69 693 -66
rect 597 -86 603 -69
rect 687 -86 693 -69
rect 597 -89 693 -86
rect 726 -69 822 -66
rect 726 -86 732 -69
rect 816 -86 822 -69
rect 726 -89 822 -86
rect 855 -69 951 -66
rect 855 -86 861 -69
rect 945 -86 951 -69
rect 855 -89 951 -86
rect 984 -69 1080 -66
rect 984 -86 990 -69
rect 1074 -86 1080 -69
rect 984 -89 1080 -86
rect 1113 -69 1209 -66
rect 1113 -86 1119 -69
rect 1203 -86 1209 -69
rect 1113 -89 1209 -86
rect 1242 -69 1338 -66
rect 1242 -86 1248 -69
rect 1332 -86 1338 -69
rect 1242 -89 1338 -86
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 21 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
