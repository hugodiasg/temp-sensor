magic
tech sky130A
magscale 1 2
timestamp 1675569099
<< metal4 >>
rect -8407 7399 -3069 7440
rect -8407 2681 -3325 7399
rect -3089 2681 -3069 7399
rect -8407 2640 -3069 2681
rect -2669 7399 2669 7440
rect -2669 2681 2413 7399
rect 2649 2681 2669 7399
rect -2669 2640 2669 2681
rect 3069 7399 8407 7440
rect 3069 2681 8151 7399
rect 8387 2681 8407 7399
rect 3069 2640 8407 2681
rect -8407 2359 -3069 2400
rect -8407 -2359 -3325 2359
rect -3089 -2359 -3069 2359
rect -8407 -2400 -3069 -2359
rect -2669 2359 2669 2400
rect -2669 -2359 2413 2359
rect 2649 -2359 2669 2359
rect -2669 -2400 2669 -2359
rect 3069 2359 8407 2400
rect 3069 -2359 8151 2359
rect 8387 -2359 8407 2359
rect 3069 -2400 8407 -2359
rect -8407 -2681 -3069 -2640
rect -8407 -7399 -3325 -2681
rect -3089 -7399 -3069 -2681
rect -8407 -7440 -3069 -7399
rect -2669 -2681 2669 -2640
rect -2669 -7399 2413 -2681
rect 2649 -7399 2669 -2681
rect -2669 -7440 2669 -7399
rect 3069 -2681 8407 -2640
rect 3069 -7399 8151 -2681
rect 8387 -7399 8407 -2681
rect 3069 -7440 8407 -7399
<< via4 >>
rect -3325 2681 -3089 7399
rect 2413 2681 2649 7399
rect 8151 2681 8387 7399
rect -3325 -2359 -3089 2359
rect 2413 -2359 2649 2359
rect 8151 -2359 8387 2359
rect -3325 -7399 -3089 -2681
rect 2413 -7399 2649 -2681
rect 8151 -7399 8387 -2681
<< mimcap2 >>
rect -8327 7320 -3687 7360
rect -8327 2760 -8287 7320
rect -3727 2760 -3687 7320
rect -8327 2720 -3687 2760
rect -2589 7320 2051 7360
rect -2589 2760 -2549 7320
rect 2011 2760 2051 7320
rect -2589 2720 2051 2760
rect 3149 7320 7789 7360
rect 3149 2760 3189 7320
rect 7749 2760 7789 7320
rect 3149 2720 7789 2760
rect -8327 2280 -3687 2320
rect -8327 -2280 -8287 2280
rect -3727 -2280 -3687 2280
rect -8327 -2320 -3687 -2280
rect -2589 2280 2051 2320
rect -2589 -2280 -2549 2280
rect 2011 -2280 2051 2280
rect -2589 -2320 2051 -2280
rect 3149 2280 7789 2320
rect 3149 -2280 3189 2280
rect 7749 -2280 7789 2280
rect 3149 -2320 7789 -2280
rect -8327 -2760 -3687 -2720
rect -8327 -7320 -8287 -2760
rect -3727 -7320 -3687 -2760
rect -8327 -7360 -3687 -7320
rect -2589 -2760 2051 -2720
rect -2589 -7320 -2549 -2760
rect 2011 -7320 2051 -2760
rect -2589 -7360 2051 -7320
rect 3149 -2760 7789 -2720
rect 3149 -7320 3189 -2760
rect 7749 -7320 7789 -2760
rect 3149 -7360 7789 -7320
<< mimcap2contact >>
rect -8287 2760 -3727 7320
rect -2549 2760 2011 7320
rect 3189 2760 7749 7320
rect -8287 -2280 -3727 2280
rect -2549 -2280 2011 2280
rect 3189 -2280 7749 2280
rect -8287 -7320 -3727 -2760
rect -2549 -7320 2011 -2760
rect 3189 -7320 7749 -2760
<< metal5 >>
rect -6167 7344 -5847 7560
rect -3367 7399 -3047 7560
rect -8311 7320 -3703 7344
rect -8311 2760 -8287 7320
rect -3727 2760 -3703 7320
rect -8311 2736 -3703 2760
rect -6167 2304 -5847 2736
rect -3367 2681 -3325 7399
rect -3089 2681 -3047 7399
rect -429 7344 -109 7560
rect 2371 7399 2691 7560
rect -2573 7320 2035 7344
rect -2573 2760 -2549 7320
rect 2011 2760 2035 7320
rect -2573 2736 2035 2760
rect -3367 2359 -3047 2681
rect -8311 2280 -3703 2304
rect -8311 -2280 -8287 2280
rect -3727 -2280 -3703 2280
rect -8311 -2304 -3703 -2280
rect -6167 -2736 -5847 -2304
rect -3367 -2359 -3325 2359
rect -3089 -2359 -3047 2359
rect -429 2304 -109 2736
rect 2371 2681 2413 7399
rect 2649 2681 2691 7399
rect 5309 7344 5629 7560
rect 8109 7399 8429 7560
rect 3165 7320 7773 7344
rect 3165 2760 3189 7320
rect 7749 2760 7773 7320
rect 3165 2736 7773 2760
rect 2371 2359 2691 2681
rect -2573 2280 2035 2304
rect -2573 -2280 -2549 2280
rect 2011 -2280 2035 2280
rect -2573 -2304 2035 -2280
rect -3367 -2681 -3047 -2359
rect -8311 -2760 -3703 -2736
rect -8311 -7320 -8287 -2760
rect -3727 -7320 -3703 -2760
rect -8311 -7344 -3703 -7320
rect -6167 -7560 -5847 -7344
rect -3367 -7399 -3325 -2681
rect -3089 -7399 -3047 -2681
rect -429 -2736 -109 -2304
rect 2371 -2359 2413 2359
rect 2649 -2359 2691 2359
rect 5309 2304 5629 2736
rect 8109 2681 8151 7399
rect 8387 2681 8429 7399
rect 8109 2359 8429 2681
rect 3165 2280 7773 2304
rect 3165 -2280 3189 2280
rect 7749 -2280 7773 2280
rect 3165 -2304 7773 -2280
rect 2371 -2681 2691 -2359
rect -2573 -2760 2035 -2736
rect -2573 -7320 -2549 -2760
rect 2011 -7320 2035 -2760
rect -2573 -7344 2035 -7320
rect -3367 -7560 -3047 -7399
rect -429 -7560 -109 -7344
rect 2371 -7399 2413 -2681
rect 2649 -7399 2691 -2681
rect 5309 -2736 5629 -2304
rect 8109 -2359 8151 2359
rect 8387 -2359 8429 2359
rect 8109 -2681 8429 -2359
rect 3165 -2760 7773 -2736
rect 3165 -7320 3189 -2760
rect 7749 -7320 7773 -2760
rect 3165 -7344 7773 -7320
rect 2371 -7560 2691 -7399
rect 5309 -7560 5629 -7344
rect 8109 -7399 8151 -2681
rect 8387 -7399 8429 -2681
rect 8109 -7560 8429 -7399
<< properties >>
string FIXED_BBOX 3069 2640 7869 7440
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.2 l 23.2 val 1.094k carea 2.00 cperi 0.19 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
