magic
tech sky130A
magscale 1 2
timestamp 1643995138
<< metal4 >>
rect 12800 -2000 14800 9800
<< metal5 >>
rect 0 20600 22600 22600
rect 0 18000 20000 20000
rect 0 2000 2000 18000
rect 2600 15400 17400 17400
rect 2600 4600 4600 15400
rect 5200 12800 14800 14800
rect 5200 7200 7200 12800
rect 12800 7800 14800 12800
rect 15400 7200 17400 15400
rect 5200 5200 17400 7200
rect 18000 4600 20000 18000
rect 2600 2600 20000 4600
rect 20600 2000 22600 20600
rect 0 0 22600 2000
<< labels >>
flabel metal5 746 21555 756 21585 0 FreeSans 1600 0 0 0 p1
port 0 nsew
flabel metal4 13753 -1378 13753 -1378 0 FreeSans 1600 0 0 0 p2
port 1 nsew
<< properties >>
string device l0
<< end >>
