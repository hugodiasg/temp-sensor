** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer_tb-ac.sch
**.subckt impedance-transformer_tb-ac
Vin1 net1 GND DC 0 AC 1
R3 ns12 GND 50 m=1
R4 ns22 net1 50 m=1
x1 ns11 ns12 GND impedance-transformer
x2 ns21 ns22 GND impedance-transformer
R1 net2 ns11 172.2 m=1
R2 GND ns21 172.2 m=1
Vin2 net2 GND DC 0 AC 1
**** begin user architecture code



.ac lin 1MEG 1.5G 4G
.control
destroy all
set units=degrees
run

set color0=white
set color1=black

let z0=50
let zl=169

* Find two S parameters from test circuit
let s11 = v(ns11)
let s12 = v(ns12)
let s21 = v(ns21)
let s22 = v(ns22)

* Extract Y parameters
*let StoYDelS = ((1+s11)*(1+s22)-s12*s21)*z0
*let y11 = ((1+s22)*(1-s11)+s12*s21/StoYDelS
*let y12=-2*s12/StoYDelS
*let y21=-2*s21/StoYDelS
*let y22 = ((1+s11)*(1-s22)+s12+s21)/StoYDelS

* Extract Z parameters
let StoZDelS = ((1-s11)*(1-s22)-s12*s21)/z0
let z11 = ((1+s11)*(1-s22)+s12*s21)/StoZDelS
let z12 = 2*s12/StoZDelS
let z21 = 2*s21/StoZDelS
let z22=((1-s11)*(1+s22)+s12*s21)/StoZDelS

*plot z11
*plot z12
*plot z21
*plot z22 xlimit 2.4G 2.5G
*plot ph(z22) xlimit 2.4G 2.5G
*plot z22
*plot smith z22
let z_in =z11-z12*z21/(z22+z0)
plot ph(z_in)
plot mag(z_in)
let z_output=z22-(z12*z21/(z11+zl))
plot ph(z_output)
plot mag(z_output)
let gamma=(mag(z_output)-mag(z_in))/(mag(z_output)+mag(z_in))
plot gamma*100
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer.sym # of pins=3
** sym_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer.sym
** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer.sch
.subckt impedance-transformer  in out gnd
*.iopin gnd
*.iopin in
*.iopin out
XC0 in gnd sky130_fd_pr__cap_mim_m3_2 W=24.43 L=24.43 MF=9 m=9
XC1 out gnd sky130_fd_pr__cap_mim_m3_2 W=24.962 L=24.962 MF=16 m=16
x1 in out l1
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sym
*+ # of pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sch
.subckt l1  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 592.7p m=1
Cs1 p1 net1 26.83f m=1
Cs2 p2 net2 24.25f m=1
Rs1 net1 GND 65.02 m=1
Rs2 net2 GND 14.4 m=1
R1 p2 net3 2.935 m=1
.ends

.GLOBAL GND
.end
