magic
tech sky130A
magscale 1 2
timestamp 1668740706
<< pwell >>
rect -425 -660 425 660
<< nmos >>
rect -229 -450 -29 450
rect 29 -450 229 450
<< ndiff >>
rect -287 438 -229 450
rect -287 -438 -275 438
rect -241 -438 -229 438
rect -287 -450 -229 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 229 438 287 450
rect 229 -438 241 438
rect 275 -438 287 438
rect 229 -450 287 -438
<< ndiffc >>
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
<< psubdiff >>
rect -389 590 -293 624
rect 293 590 389 624
rect -389 528 -355 590
rect 355 528 389 590
rect -389 -590 -355 -528
rect 355 -590 389 -528
rect -389 -624 -293 -590
rect 293 -624 389 -590
<< psubdiffcont >>
rect -293 590 293 624
rect -389 -528 -355 528
rect 355 -528 389 528
rect -293 -624 293 -590
<< poly >>
rect -229 522 -29 538
rect -229 488 -213 522
rect -45 488 -29 522
rect -229 450 -29 488
rect 29 522 229 538
rect 29 488 45 522
rect 213 488 229 522
rect 29 450 229 488
rect -229 -488 -29 -450
rect -229 -522 -213 -488
rect -45 -522 -29 -488
rect -229 -538 -29 -522
rect 29 -488 229 -450
rect 29 -522 45 -488
rect 213 -522 229 -488
rect 29 -538 229 -522
<< polycont >>
rect -213 488 -45 522
rect 45 488 213 522
rect -213 -522 -45 -488
rect 45 -522 213 -488
<< locali >>
rect -389 590 -293 624
rect 293 590 389 624
rect -389 528 -355 590
rect 355 528 389 590
rect -229 488 -213 522
rect -45 488 -29 522
rect 29 488 45 522
rect 213 488 229 522
rect -275 438 -241 454
rect -275 -454 -241 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 241 438 275 454
rect 241 -454 275 -438
rect -229 -522 -213 -488
rect -45 -522 -29 -488
rect 29 -522 45 -488
rect 213 -522 229 -488
rect -389 -590 -355 -528
rect 355 -590 389 -528
rect -389 -624 -293 -590
rect 293 -624 389 -590
<< viali >>
rect -213 488 -45 522
rect 45 488 213 522
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
rect -213 -522 -45 -488
rect 45 -522 213 -488
<< metal1 >>
rect -225 522 -33 528
rect -225 488 -213 522
rect -45 488 -33 522
rect -225 482 -33 488
rect 33 522 225 528
rect 33 488 45 522
rect 213 488 225 522
rect 33 482 225 488
rect -281 438 -235 450
rect -281 -438 -275 438
rect -241 -438 -235 438
rect -281 -450 -235 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 235 438 281 450
rect 235 -438 241 438
rect 275 -438 281 438
rect 235 -450 281 -438
rect -225 -488 -33 -482
rect -225 -522 -213 -488
rect -45 -522 -33 -488
rect -225 -528 -33 -522
rect 33 -488 225 -482
rect 33 -522 45 -488
rect 213 -522 225 -488
rect 33 -528 225 -522
<< properties >>
string FIXED_BBOX -372 -607 372 607
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.5 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
