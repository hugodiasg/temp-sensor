* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[10] io_analog[3]
+ io_analog[7] io_analog[8] io_analog[9] io_analog[5] io_analog[6] io_clamp_high[0]
+ io_clamp_high[1] io_clamp_high[2] io_clamp_low[0] io_clamp_low[1] io_clamp_low[2]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26]
+ io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0]
+ io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[14] io_in_3v3[15]
+ io_in_3v3[16] io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1] io_in_3v3[20]
+ io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25] io_in_3v3[26]
+ io_in_3v3[2] io_in_3v3[3] io_in_3v3[4] io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8]
+ io_in_3v3[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0]
+ la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2
+ user_irq[0] user_irq[1] user_irq[2] vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i io_analog[1] io_in[13]
+ io_analog[0] io_analog[2] io_analog[4] vccd1
X0 a_448090_652460# a_448256_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X1 device-complete_0.buffer_0.b device-complete_0.buffer_0.b vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 io_analog[0] a_449985_647995# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 a_449355_647995# a_448165_647995# a_449246_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=21.2 ps=177 w=1 l=1
X5 a_448789_648361# vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X6 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=1
X7 a_448777_647995# a_448331_647995# a_448681_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X8 io_analog[4] device-complete_0.vtd device-complete_0.vtd io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_449408_648361# a_448331_647995# a_449246_647995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.a vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X12 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.a vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X13 vdda1 device-complete_0.buffer_0.a device-complete_0.buffer_0.a vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a_450228_652460# a_450394_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X15 io_analog[4] io_analog[4] io_analog[4] io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=5.22 ps=41.2 w=2 l=1
X16 io_analog[1] device-complete_0.buffer_0.b vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X17 vdda1 device-complete_0.buffer_0.b device-complete_0.buffer_0.b vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 vccd1 a_449421_647969# a_449985_647995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X19 device-complete_0.vtd device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X20 a_448306_650292# a_448472_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X21 device-complete_0.sensor_0.c device-complete_0.sensor_0.c device-complete_0.sensor_0.c vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=1
X22 vssa1 io_analog[2] io_analog[2] vssa1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 vssa1 vccd1 a_448943_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_448090_652460# io_analog[1] vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X25 vdda1 device-complete_0.sensor_0.a device-complete_0.sensor_0.a vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X26 device-complete_0.buffer_0.d device-complete_0.buffer_0.d device-complete_0.buffer_0.d vdda1 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=17.4 ps=122 w=15 l=1
X27 vccd1 a_449246_647995# a_449421_647969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 device-complete_0.sensor_0.a device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X29 device-complete_0.sensor_0.a device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X30 a_450560_652460# device-complete_0.sigma-delta_0.x1.Q vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X31 io_analog[4] io_analog[4] io_analog[4] io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X32 device-complete_0.vtd device-complete_0.vtd io_analog[4] io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_448638_650292# a_448804_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X34 a_449086_652460# device-complete_0.sigma-delta_0.in_int vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X35 a_448422_652460# a_448588_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X36 a_448899_648237# a_448681_647995# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X37 device-complete_0.sensor_0.c device-complete_0.sensor_0.a device-complete_0.sensor_0.d vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X38 device-complete_0.buffer_0.a device-complete_0.buffer_0.a device-complete_0.buffer_0.a vssa1 sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0.96 ps=7.28 w=1.5 l=0.15
X39 a_448422_652460# a_448256_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X40 vccd1 io_in[13] a_448165_647995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X41 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X42 device-complete_0.buffer_0.a device-complete_0.buffer_0.a vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X43 io_analog[2] io_analog[2] io_analog[2] vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.58 ps=5.16 w=1 l=1
X44 a_448586_647995# device-complete_0.sigma-delta_0.x1.D vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X45 a_448943_647995# a_448899_648237# a_448777_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X46 vssa1 device-complete_0.buffer_0.d io_analog[1] vssa1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 device-complete_0.sensor_0.b device-complete_0.vtd device-complete_0.sensor_0.c vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X48 io_analog[4] device-complete_0.vtd device-complete_0.vtd io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X49 device-complete_0.buffer_0.d device-complete_0.buffer_0.d device-complete_0.buffer_0.d vdda1 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0 w=15 l=1
X50 vssa1 a_449421_647969# a_449985_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X51 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.a vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X52 a_450560_652460# a_450394_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X53 vdda1 vdda1 vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=17.1 ps=130 w=1 l=1
X54 io_analog[1] io_analog[1] io_analog[1] vdda1 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=17.4 ps=122 w=15 l=1
X55 device-complete_0.sigma-delta_0.in_int vssa1 sky130_fd_pr__cap_mim_m3_2 l=27.2 w=27.2
X56 vccd1 a_448899_648237# a_448789_648361# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X57 vdda1 io_analog[3] sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X58 vdda1 device-complete_0.buffer_0.b device-complete_0.buffer_0.b vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X59 vdda1 a_439666_676526# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=5
X60 a_449246_647995# a_448165_647995# a_448899_648237# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X61 vssa1 device-complete_0.sensor_0.b device-complete_0.vtd vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X62 device-complete_0.vtd device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X63 vssa1 device-complete_0.sensor_0.b device-complete_0.vtd vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X64 device-complete_0.buffer_0.b device-complete_0.buffer_0.b device-complete_0.buffer_0.b vssa1 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.96 ps=7.28 w=1.5 l=0.15
X65 a_448754_652460# a_448588_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X66 device-complete_0.sensor_0.c device-complete_0.vtd device-complete_0.sensor_0.b vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X67 device-complete_0.sensor_0.a device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X68 vdda1 device-complete_0.vtd io_analog[4] vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X69 vssa1 io_in[13] a_448165_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X70 a_448681_647995# a_448165_647995# a_448586_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X71 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X72 a_448970_650292# a_448804_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X73 device-complete_0.buffer_0.d device-complete_0.buffer_0.a vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X74 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X75 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X76 vssa1 device-complete_0.buffer_0.d device-complete_0.buffer_0.d vssa1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X77 device-complete_0.vtd device-complete_0.vtd io_analog[4] io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X78 io_analog[0] a_449985_647995# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X79 a_449564_652460# device-complete_0.sigma-delta_0.in_int vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X80 device-complete_0.buffer_0.a device-complete_0.buffer_0.a vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X81 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.a vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X82 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X83 vdda1 device-complete_0.buffer_0.b io_analog[1] vdda1 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X84 a_449421_647969# a_449246_647995# a_449600_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X85 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X86 device-complete_0.buffer_0.b device-complete_0.buffer_0.b device-complete_0.buffer_0.b vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=1.16 ps=10.3 w=1 l=1
X87 a_448754_652460# a_448920_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X88 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X89 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X90 vssa1 io_analog[0] io_analog[3] vssa1 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X91 device-complete_0.sensor_0.b device-complete_0.vtd device-complete_0.sensor_0.c vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X92 vccd1 a_449421_647969# a_449408_648361# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X93 vssa1 device-complete_0.sensor_0.b device-complete_0.vtd vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X94 device-complete_0.buffer_0.d device-complete_0.buffer_0.d vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 io_analog[4] device-complete_0.vtd device-complete_0.vtd io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X96 vdda1 vdda1 vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X97 vdda1 io_analog[3] sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X98 device-complete_0.sensor_0.d device-complete_0.sensor_0.a device-complete_0.sensor_0.c vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X99 device-complete_0.sensor_0.a device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X100 device-complete_0.sensor_0.d device-complete_0.sensor_0.a device-complete_0.sensor_0.c vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X101 a_448899_648237# a_448681_647995# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X102 vdda1 vdda1 vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X103 vssa1 device-complete_0.sigma-delta_0.in_comp device-complete_0.sigma-delta_0.x1.D vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X104 a_449896_652460# a_449730_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X105 io_analog[1] device-complete_0.buffer_0.d vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_448789_648361# a_448165_647995# a_448681_647995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X107 device-complete_0.sensor_0.c device-complete_0.vtd device-complete_0.sensor_0.b vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X108 vdda1 io_analog[3] sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X109 a_449600_647995# vccd1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X110 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X111 a_449564_652460# a_449730_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X112 a_448331_647995# a_448165_647995# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X113 io_analog[4] device-complete_0.vtd device-complete_0.vtd io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X114 device-complete_0.sigma-delta_0.x1.Q a_449421_647969# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X115 vdda1 device-complete_0.buffer_0.a device-complete_0.buffer_0.a vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X116 device-complete_0.buffer_0.b io_analog[4] device-complete_0.buffer_0.c vssa1 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X117 io_analog[1] io_analog[1] io_analog[1] vdda1 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0 w=15 l=1
X118 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X119 a_448970_650292# a_449136_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X120 device-complete_0.sigma-delta_0.x1.Q a_449421_647969# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.213 ps=1.67 w=1 l=0.15
X121 a_450228_652460# a_450062_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X122 vdda1 device-complete_0.buffer_0.b device-complete_0.buffer_0.b vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X123 vdda1 vdda1 vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X124 device-complete_0.buffer_0.c device-complete_0.buffer_0.c device-complete_0.buffer_0.c vssa1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=1.08 ps=8.82 w=1 l=1
X125 a_448306_650292# a_448140_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X126 device-complete_0.buffer_0.c io_analog[1] device-complete_0.buffer_0.a vssa1 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X127 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X128 vssa1 vssa1 vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=1
X129 a_448681_647995# a_448331_647995# a_448586_647995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X130 vssa1 device-complete_0.sensor_0.b device-complete_0.vtd vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X131 device-complete_0.vtd device-complete_0.vtd io_analog[4] io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X132 device-complete_0.sensor_0.c device-complete_0.sensor_0.a device-complete_0.sensor_0.d vdda1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X133 device-complete_0.buffer_0.a device-complete_0.buffer_0.a device-complete_0.buffer_0.a vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=1.16 ps=10.3 w=1 l=1
X134 vdda1 vdda1 vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X135 a_449246_647995# a_448331_647995# a_448899_648237# vssa1 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X136 device-complete_0.vtd device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X137 device-complete_0.vtd device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X138 device-complete_0.sensor_0.d device-complete_0.vtd vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X139 device-complete_0.buffer_0.b device-complete_0.buffer_0.b vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X140 device-complete_0.buffer_0.c io_analog[2] vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X141 a_448586_647995# device-complete_0.sigma-delta_0.x1.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X142 vdda1 device-complete_0.sigma-delta_0.in_comp device-complete_0.sigma-delta_0.x1.D vdda1 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X143 device-complete_0.sensor_0.a device-complete_0.sensor_0.a vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X144 a_449896_652460# a_450062_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X145 vdda1 device-complete_0.buffer_0.a device-complete_0.buffer_0.d vdda1 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X146 io_analog[1] device-complete_0.buffer_0.d sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X147 device-complete_0.sigma-delta_0.in_int a_448140_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X148 device-complete_0.vtd device-complete_0.vtd io_analog[4] io_analog[4] sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X149 device-complete_0.sigma-delta_0.in_comp vssa1 sky130_fd_pr__cap_mim_m3_2 l=27.2 w=27.2
X150 vssa1 a_449421_647969# a_449355_647995# vssa1 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X151 a_449421_647969# vccd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X152 a_448331_647995# a_448165_647995# vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X153 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X154 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X155 device-complete_0.sigma-delta_0.in_comp a_449136_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X156 a_448638_650292# a_448472_649460# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=2
X157 a_449086_652460# a_448920_651128# vssa1 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X158 device-complete_0.buffer_0.a device-complete_0.buffer_0.a vdda1 vdda1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X159 vssa1 device-complete_0.sensor_0.b device-complete_0.sensor_0.b vssa1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

