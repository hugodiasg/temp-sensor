magic
tech sky130A
magscale 1 2
timestamp 1645799662
<< metal4 >>
rect -2379 9309 2379 9350
rect -2379 4791 2123 9309
rect 2359 4791 2379 9309
rect -2379 4750 2379 4791
rect -2379 4609 2379 4650
rect -2379 91 2123 4609
rect 2359 91 2379 4609
rect -2379 50 2379 91
rect -2379 -91 2379 -50
rect -2379 -4609 2123 -91
rect 2359 -4609 2379 -91
rect -2379 -4650 2379 -4609
rect -2379 -4791 2379 -4750
rect -2379 -9309 2123 -4791
rect 2359 -9309 2379 -4791
rect -2379 -9350 2379 -9309
<< via4 >>
rect 2123 4791 2359 9309
rect 2123 91 2359 4609
rect 2123 -4609 2359 -91
rect 2123 -9309 2359 -4791
<< mimcap2 >>
rect -2279 9210 2121 9250
rect -2279 4890 -1807 9210
rect 1649 4890 2121 9210
rect -2279 4850 2121 4890
rect -2279 4510 2121 4550
rect -2279 190 -1807 4510
rect 1649 190 2121 4510
rect -2279 150 2121 190
rect -2279 -190 2121 -150
rect -2279 -4510 -1807 -190
rect 1649 -4510 2121 -190
rect -2279 -4550 2121 -4510
rect -2279 -4890 2121 -4850
rect -2279 -9210 -1807 -4890
rect 1649 -9210 2121 -4890
rect -2279 -9250 2121 -9210
<< mimcap2contact >>
rect -1807 4890 1649 9210
rect -1807 190 1649 4510
rect -1807 -4510 1649 -190
rect -1807 -9210 1649 -4890
<< metal5 >>
rect -239 9234 81 9400
rect 2081 9309 2401 9400
rect -1831 9210 1673 9234
rect -1831 4890 -1807 9210
rect 1649 4890 1673 9210
rect -1831 4866 1673 4890
rect -239 4534 81 4866
rect 2081 4791 2123 9309
rect 2359 4791 2401 9309
rect 2081 4609 2401 4791
rect -1831 4510 1673 4534
rect -1831 190 -1807 4510
rect 1649 190 1673 4510
rect -1831 166 1673 190
rect -239 -166 81 166
rect 2081 91 2123 4609
rect 2359 91 2401 4609
rect 2081 -91 2401 91
rect -1831 -190 1673 -166
rect -1831 -4510 -1807 -190
rect 1649 -4510 1673 -190
rect -1831 -4534 1673 -4510
rect -239 -4866 81 -4534
rect 2081 -4609 2123 -91
rect 2359 -4609 2401 -91
rect 2081 -4791 2401 -4609
rect -1831 -4890 1673 -4866
rect -1831 -9210 -1807 -4890
rect 1649 -9210 1673 -4890
rect -1831 -9234 1673 -9210
rect -239 -9400 81 -9234
rect 2081 -9309 2123 -4791
rect 2359 -9309 2401 -4791
rect 2081 -9400 2401 -9309
<< properties >>
string FIXED_BBOX -2379 4750 2221 9350
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
