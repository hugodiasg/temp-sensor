magic
tech sky130A
magscale 1 2
timestamp 1646064585
<< metal4 >>
rect -2757 10821 2757 10862
rect -2757 5547 2501 10821
rect 2737 5547 2757 10821
rect -2757 5506 2757 5547
rect -2757 5365 2757 5406
rect -2757 91 2501 5365
rect 2737 91 2757 5365
rect -2757 50 2757 91
rect -2757 -91 2757 -50
rect -2757 -5365 2501 -91
rect 2737 -5365 2757 -91
rect -2757 -5406 2757 -5365
rect -2757 -5547 2757 -5506
rect -2757 -10821 2501 -5547
rect 2737 -10821 2757 -5547
rect -2757 -10862 2757 -10821
<< via4 >>
rect 2501 5547 2737 10821
rect 2501 91 2737 5365
rect 2501 -5365 2737 -91
rect 2501 -10821 2737 -5547
<< mimcap2 >>
rect -2657 10722 2499 10762
rect -2657 5646 -2109 10722
rect 1951 5646 2499 10722
rect -2657 5606 2499 5646
rect -2657 5266 2499 5306
rect -2657 190 -2109 5266
rect 1951 190 2499 5266
rect -2657 150 2499 190
rect -2657 -190 2499 -150
rect -2657 -5266 -2109 -190
rect 1951 -5266 2499 -190
rect -2657 -5306 2499 -5266
rect -2657 -5646 2499 -5606
rect -2657 -10722 -2109 -5646
rect 1951 -10722 2499 -5646
rect -2657 -10762 2499 -10722
<< mimcap2contact >>
rect -2109 5646 1951 10722
rect -2109 190 1951 5266
rect -2109 -5266 1951 -190
rect -2109 -10722 1951 -5646
<< metal5 >>
rect -239 10746 81 10912
rect 2459 10821 2779 10912
rect -2133 10722 1975 10746
rect -2133 5646 -2109 10722
rect 1951 5646 1975 10722
rect -2133 5622 1975 5646
rect -239 5290 81 5622
rect 2459 5547 2501 10821
rect 2737 5547 2779 10821
rect 2459 5365 2779 5547
rect -2133 5266 1975 5290
rect -2133 190 -2109 5266
rect 1951 190 1975 5266
rect -2133 166 1975 190
rect -239 -166 81 166
rect 2459 91 2501 5365
rect 2737 91 2779 5365
rect 2459 -91 2779 91
rect -2133 -190 1975 -166
rect -2133 -5266 -2109 -190
rect 1951 -5266 1975 -190
rect -2133 -5290 1975 -5266
rect -239 -5622 81 -5290
rect 2459 -5365 2501 -91
rect 2737 -5365 2779 -91
rect 2459 -5547 2779 -5365
rect -2133 -5646 1975 -5622
rect -2133 -10722 -2109 -5646
rect 1951 -10722 1975 -5646
rect -2133 -10746 1975 -10722
rect -239 -10912 81 -10746
rect 2459 -10821 2501 -5547
rect 2737 -10821 2779 -5547
rect 2459 -10912 2779 -10821
<< properties >>
string FIXED_BBOX -2757 5506 2599 10862
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.781 l 25.781 val 1.348k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
