magic
tech sky130A
magscale 1 2
timestamp 1646183319
<< metal4 >>
rect -2590 10153 2590 10194
rect -2590 5213 2334 10153
rect 2570 5213 2590 10153
rect -2590 5172 2590 5213
rect -2590 5031 2590 5072
rect -2590 91 2334 5031
rect 2570 91 2590 5031
rect -2590 50 2590 91
rect -2590 -91 2590 -50
rect -2590 -5031 2334 -91
rect 2570 -5031 2590 -91
rect -2590 -5072 2590 -5031
rect -2590 -5213 2590 -5172
rect -2590 -10153 2334 -5213
rect 2570 -10153 2590 -5213
rect -2590 -10194 2590 -10153
<< via4 >>
rect 2334 5213 2570 10153
rect 2334 91 2570 5031
rect 2334 -5031 2570 -91
rect 2334 -10153 2570 -5213
<< mimcap2 >>
rect -2490 10054 2332 10094
rect -2490 5312 -1976 10054
rect 1818 5312 2332 10054
rect -2490 5272 2332 5312
rect -2490 4932 2332 4972
rect -2490 190 -1976 4932
rect 1818 190 2332 4932
rect -2490 150 2332 190
rect -2490 -190 2332 -150
rect -2490 -4932 -1976 -190
rect 1818 -4932 2332 -190
rect -2490 -4972 2332 -4932
rect -2490 -5312 2332 -5272
rect -2490 -10054 -1976 -5312
rect 1818 -10054 2332 -5312
rect -2490 -10094 2332 -10054
<< mimcap2contact >>
rect -1976 5312 1818 10054
rect -1976 190 1818 4932
rect -1976 -4932 1818 -190
rect -1976 -10054 1818 -5312
<< metal5 >>
rect -239 10078 81 10244
rect 2292 10153 2612 10244
rect -2000 10054 1842 10078
rect -2000 5312 -1976 10054
rect 1818 5312 1842 10054
rect -2000 5288 1842 5312
rect -239 4956 81 5288
rect 2292 5213 2334 10153
rect 2570 5213 2612 10153
rect 2292 5031 2612 5213
rect -2000 4932 1842 4956
rect -2000 190 -1976 4932
rect 1818 190 1842 4932
rect -2000 166 1842 190
rect -239 -166 81 166
rect 2292 91 2334 5031
rect 2570 91 2612 5031
rect 2292 -91 2612 91
rect -2000 -190 1842 -166
rect -2000 -4932 -1976 -190
rect 1818 -4932 1842 -190
rect -2000 -4956 1842 -4932
rect -239 -5288 81 -4956
rect 2292 -5031 2334 -91
rect 2570 -5031 2612 -91
rect 2292 -5213 2612 -5031
rect -2000 -5312 1842 -5288
rect -2000 -10054 -1976 -5312
rect 1818 -10054 1842 -5312
rect -2000 -10078 1842 -10054
rect -239 -10244 81 -10078
rect 2292 -10153 2334 -5213
rect 2570 -10153 2612 -5213
rect 2292 -10244 2612 -10153
<< properties >>
string FIXED_BBOX -2590 5172 2432 10194
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.111 l 24.111 val 1.181k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
