magic
tech sky130A
magscale 1 2
timestamp 1656875000
<< metal3 >>
rect -2250 2172 2249 2200
rect -2250 -2172 2165 2172
rect 2229 -2172 2249 2172
rect -2250 -2200 2249 -2172
<< via3 >>
rect 2165 -2172 2229 2172
<< mimcap >>
rect -2150 2060 2050 2100
rect -2150 -2060 -2110 2060
rect 2010 -2060 2050 2060
rect -2150 -2100 2050 -2060
<< mimcapcontact >>
rect -2110 -2060 2010 2060
<< metal4 >>
rect 2149 2172 2245 2188
rect -2111 2060 2011 2061
rect -2111 -2060 -2110 2060
rect 2010 -2060 2011 2060
rect -2111 -2061 2011 -2060
rect 2149 -2172 2165 2172
rect 2229 -2172 2245 2172
rect 2149 -2188 2245 -2172
<< properties >>
string FIXED_BBOX -2250 -2200 2150 2200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 21.0 l 21.0 val 897.96 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
