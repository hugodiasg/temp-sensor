magic
tech sky130A
magscale 1 2
timestamp 1646100680
<< metal4 >>
rect -2504 7334 2504 7375
rect -2504 2566 2248 7334
rect 2484 2566 2504 7334
rect -2504 2525 2504 2566
rect -2504 2384 2504 2425
rect -2504 -2384 2248 2384
rect 2484 -2384 2504 2384
rect -2504 -2425 2504 -2384
rect -2504 -2566 2504 -2525
rect -2504 -7334 2248 -2566
rect 2484 -7334 2504 -2566
rect -2504 -7375 2504 -7334
<< via4 >>
rect 2248 2566 2484 7334
rect 2248 -2384 2484 2384
rect 2248 -7334 2484 -2566
<< mimcap2 >>
rect -2404 7235 2246 7275
rect -2404 2665 -1907 7235
rect 1749 2665 2246 7235
rect -2404 2625 2246 2665
rect -2404 2285 2246 2325
rect -2404 -2285 -1907 2285
rect 1749 -2285 2246 2285
rect -2404 -2325 2246 -2285
rect -2404 -2665 2246 -2625
rect -2404 -7235 -1907 -2665
rect 1749 -7235 2246 -2665
rect -2404 -7275 2246 -7235
<< mimcap2contact >>
rect -1907 2665 1749 7235
rect -1907 -2285 1749 2285
rect -1907 -7235 1749 -2665
<< metal5 >>
rect -239 7259 81 7425
rect 2206 7334 2526 7425
rect -1931 7235 1773 7259
rect -1931 2665 -1907 7235
rect 1749 2665 1773 7235
rect -1931 2641 1773 2665
rect -239 2309 81 2641
rect 2206 2566 2248 7334
rect 2484 2566 2526 7334
rect 2206 2384 2526 2566
rect -1931 2285 1773 2309
rect -1931 -2285 -1907 2285
rect 1749 -2285 1773 2285
rect -1931 -2309 1773 -2285
rect -239 -2641 81 -2309
rect 2206 -2384 2248 2384
rect 2484 -2384 2526 2384
rect 2206 -2566 2526 -2384
rect -1931 -2665 1773 -2641
rect -1931 -7235 -1907 -2665
rect 1749 -7235 1773 -2665
rect -1931 -7259 1773 -7235
rect -239 -7425 81 -7259
rect 2206 -7334 2248 -2566
rect 2484 -7334 2526 -2566
rect 2206 -7425 2526 -7334
<< properties >>
string FIXED_BBOX -2504 2525 2346 7375
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.252 l 23.252 val 1.098k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
