** sch_path: /foss/designs/temp-sensor/ask_modulator/xschem/ask-modulator-pex_tb-tran.sch
**.subckt ask-modulator-pex_tb-tran
Vdd vd GND 1.8
V1 in GND pulse 0 1.8 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 '
x1 vd out in GND ask-modulator-pex
**** begin user architecture code




.tran 40p 150n

.control
destroy all
run

set color0=white
set color1=black

let id =-i(vdd)
*plot id
plot in
plot out

* FFT
linearize out
fft out
plot mag(out) xlimit 1.7G 4G ylimit 0 50u
.endc

 .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/temp-sensor/ask_modulator/xschem/ask-modulator-pex.sym # of
*+ pins=4
** sym_path: /foss/designs/temp-sensor/ask_modulator/xschem/ask-modulator-pex.sym
** sch_path: /foss/designs/temp-sensor/ask_modulator/xschem/ask-modulator-pex.sch
.subckt ask-modulator-pex vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
**** begin user architecture code


* NGSPICE file created from ask-modulator.ext - technology: sky130A

*.subckt ask-modulator gnd in out vd
X0 vd.t1 out.t2 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X1 vd.t0 a_6666_12466# gnd.t0 sky130_fd_pr__res_xhigh_po_0p35 l=5
X2 vd.t2 out.t1 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X3 gnd.t2 in.t0 out.t3 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X4 vd.t3 out.t0 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
R0 vd.n2 vd.t0 9.57793
R1 vd vd.n2 0.156465
R2 vd.n0 vd.t3 0.0686501
R3 vd.n1 vd.n0 0.06865
R4 vd.n2 vd.n1 0.00834818
R5 vd.n0 vd.t1 0.000500086
R6 vd.n1 vd.t2 0.000500086
R7 out.n2 out.t3 8.96122
R8 out.n2 out.n1 1.04919
R9 out.n0 out.t1 0.506271
R10 out.n1 out.n0 0.480533
R11 out.n3 out.n2 0.130708
R12 out.n3 out 0.0755
R13 out out.n3 0.063
R14 out.n0 out.t2 0.0277714
R15 out.n1 out.t0 0.0262381
R16 gnd.n12 gnd.n11 840.21
R17 gnd.n17 gnd.n14 25.7727
R18 gnd.n20 gnd.t1 25.4863
R19 gnd.n11 gnd.t0 24.3353
R20 gnd.n8 gnd.n5 24.2558
R21 gnd.n28 gnd.n27 9.15497
R22 gnd.n29 gnd.t2 8.74711
R23 gnd.n28 gnd.n26 5.56572
R24 gnd gnd.n29 3.03327
R25 gnd.n23 gnd.n12 2.30244
R26 gnd.n23 gnd.n20 0.493774
R27 gnd.n22 gnd.n21 0.288252
R28 gnd.n23 gnd.n22 0.288252
R29 gnd.n24 gnd.n1 0.202818
R30 gnd.n1 gnd.n0 0.202363
R31 gnd.n8 gnd.n7 0.130535
R32 gnd.n3 gnd.n2 0.1305
R33 gnd.t0 gnd.n3 0.1305
R34 gnd.n7 gnd.n6 0.1305
R35 gnd.n19 gnd.n18 0.10956
R36 gnd.t1 gnd.n19 0.10956
R37 gnd.n16 gnd.n15 0.10956
R38 gnd.n17 gnd.n16 0.109082
R39 gnd.n25 gnd.n24 0.0528087
R40 gnd.n26 gnd.n25 0.0523204
R41 gnd.n14 gnd.n13 0.0264102
R42 gnd.n10 gnd.n9 0.00762598
R43 gnd.n11 gnd.n10 0.00762598
R44 gnd.n5 gnd.n4 0.00762598
R45 gnd.t1 gnd.n17 0.00197408
R46 gnd.n29 gnd.n28 0.001518
R47 gnd.t0 gnd.n8 0.00146275
R48 gnd.n24 gnd.n23 0.0010093
R49 in in.t0 393.923
C0 out a_6666_12466# 0.231f
C1 out vd 0.139p
C2 out in 0.229f
C3 vd a_6666_12466# 0.138f
*.ends



**** end user architecture code
x1 vd out l0
.ends


* expanding   symbol:  /foss/designs/temp-sensor/ask_modulator/xschem/l0.sym # of pins=2
** sym_path: /foss/designs/temp-sensor/ask_modulator/xschem/l0.sym
** sch_path: /foss/designs/temp-sensor/ask_modulator/xschem/l0.sch
.subckt l0 p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 993p m=1
Cs1 p1 net1 58.53f m=1
Cs2 p2 net2 52.93f m=1
Rs1 net1 GND 24.1 m=1
Rs2 net2 GND 22.94 m=1
R1 p2 net3 3.443 m=1
.ends

.GLOBAL GND
.end
