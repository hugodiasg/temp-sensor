magic
tech sky130A
magscale 1 2
timestamp 1661301161
<< pwell >>
rect -2747 -310 2747 310
<< nmos >>
rect -2551 -100 -2351 100
rect -2293 -100 -2093 100
rect -2035 -100 -1835 100
rect -1777 -100 -1577 100
rect -1519 -100 -1319 100
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
rect 1319 -100 1519 100
rect 1577 -100 1777 100
rect 1835 -100 2035 100
rect 2093 -100 2293 100
rect 2351 -100 2551 100
<< ndiff >>
rect -2609 88 -2551 100
rect -2609 -88 -2597 88
rect -2563 -88 -2551 88
rect -2609 -100 -2551 -88
rect -2351 88 -2293 100
rect -2351 -88 -2339 88
rect -2305 -88 -2293 88
rect -2351 -100 -2293 -88
rect -2093 88 -2035 100
rect -2093 -88 -2081 88
rect -2047 -88 -2035 88
rect -2093 -100 -2035 -88
rect -1835 88 -1777 100
rect -1835 -88 -1823 88
rect -1789 -88 -1777 88
rect -1835 -100 -1777 -88
rect -1577 88 -1519 100
rect -1577 -88 -1565 88
rect -1531 -88 -1519 88
rect -1577 -100 -1519 -88
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
rect 1519 88 1577 100
rect 1519 -88 1531 88
rect 1565 -88 1577 88
rect 1519 -100 1577 -88
rect 1777 88 1835 100
rect 1777 -88 1789 88
rect 1823 -88 1835 88
rect 1777 -100 1835 -88
rect 2035 88 2093 100
rect 2035 -88 2047 88
rect 2081 -88 2093 88
rect 2035 -100 2093 -88
rect 2293 88 2351 100
rect 2293 -88 2305 88
rect 2339 -88 2351 88
rect 2293 -100 2351 -88
rect 2551 88 2609 100
rect 2551 -88 2563 88
rect 2597 -88 2609 88
rect 2551 -100 2609 -88
<< ndiffc >>
rect -2597 -88 -2563 88
rect -2339 -88 -2305 88
rect -2081 -88 -2047 88
rect -1823 -88 -1789 88
rect -1565 -88 -1531 88
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect 1531 -88 1565 88
rect 1789 -88 1823 88
rect 2047 -88 2081 88
rect 2305 -88 2339 88
rect 2563 -88 2597 88
<< psubdiff >>
rect -2711 240 -2615 274
rect 2615 240 2711 274
rect -2711 178 -2677 240
rect 2677 178 2711 240
rect -2711 -240 -2677 -178
rect 2677 -240 2711 -178
rect -2711 -274 -2615 -240
rect 2615 -274 2711 -240
<< psubdiffcont >>
rect -2615 240 2615 274
rect -2711 -178 -2677 178
rect 2677 -178 2711 178
rect -2615 -274 2615 -240
<< poly >>
rect -2551 172 -2351 188
rect -2551 138 -2535 172
rect -2367 138 -2351 172
rect -2551 100 -2351 138
rect -2293 172 -2093 188
rect -2293 138 -2277 172
rect -2109 138 -2093 172
rect -2293 100 -2093 138
rect -2035 172 -1835 188
rect -2035 138 -2019 172
rect -1851 138 -1835 172
rect -2035 100 -1835 138
rect -1777 172 -1577 188
rect -1777 138 -1761 172
rect -1593 138 -1577 172
rect -1777 100 -1577 138
rect -1519 172 -1319 188
rect -1519 138 -1503 172
rect -1335 138 -1319 172
rect -1519 100 -1319 138
rect -1261 172 -1061 188
rect -1261 138 -1245 172
rect -1077 138 -1061 172
rect -1261 100 -1061 138
rect -1003 172 -803 188
rect -1003 138 -987 172
rect -819 138 -803 172
rect -1003 100 -803 138
rect -745 172 -545 188
rect -745 138 -729 172
rect -561 138 -545 172
rect -745 100 -545 138
rect -487 172 -287 188
rect -487 138 -471 172
rect -303 138 -287 172
rect -487 100 -287 138
rect -229 172 -29 188
rect -229 138 -213 172
rect -45 138 -29 172
rect -229 100 -29 138
rect 29 172 229 188
rect 29 138 45 172
rect 213 138 229 172
rect 29 100 229 138
rect 287 172 487 188
rect 287 138 303 172
rect 471 138 487 172
rect 287 100 487 138
rect 545 172 745 188
rect 545 138 561 172
rect 729 138 745 172
rect 545 100 745 138
rect 803 172 1003 188
rect 803 138 819 172
rect 987 138 1003 172
rect 803 100 1003 138
rect 1061 172 1261 188
rect 1061 138 1077 172
rect 1245 138 1261 172
rect 1061 100 1261 138
rect 1319 172 1519 188
rect 1319 138 1335 172
rect 1503 138 1519 172
rect 1319 100 1519 138
rect 1577 172 1777 188
rect 1577 138 1593 172
rect 1761 138 1777 172
rect 1577 100 1777 138
rect 1835 172 2035 188
rect 1835 138 1851 172
rect 2019 138 2035 172
rect 1835 100 2035 138
rect 2093 172 2293 188
rect 2093 138 2109 172
rect 2277 138 2293 172
rect 2093 100 2293 138
rect 2351 172 2551 188
rect 2351 138 2367 172
rect 2535 138 2551 172
rect 2351 100 2551 138
rect -2551 -138 -2351 -100
rect -2551 -172 -2535 -138
rect -2367 -172 -2351 -138
rect -2551 -188 -2351 -172
rect -2293 -138 -2093 -100
rect -2293 -172 -2277 -138
rect -2109 -172 -2093 -138
rect -2293 -188 -2093 -172
rect -2035 -138 -1835 -100
rect -2035 -172 -2019 -138
rect -1851 -172 -1835 -138
rect -2035 -188 -1835 -172
rect -1777 -138 -1577 -100
rect -1777 -172 -1761 -138
rect -1593 -172 -1577 -138
rect -1777 -188 -1577 -172
rect -1519 -138 -1319 -100
rect -1519 -172 -1503 -138
rect -1335 -172 -1319 -138
rect -1519 -188 -1319 -172
rect -1261 -138 -1061 -100
rect -1261 -172 -1245 -138
rect -1077 -172 -1061 -138
rect -1261 -188 -1061 -172
rect -1003 -138 -803 -100
rect -1003 -172 -987 -138
rect -819 -172 -803 -138
rect -1003 -188 -803 -172
rect -745 -138 -545 -100
rect -745 -172 -729 -138
rect -561 -172 -545 -138
rect -745 -188 -545 -172
rect -487 -138 -287 -100
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -487 -188 -287 -172
rect -229 -138 -29 -100
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect -229 -188 -29 -172
rect 29 -138 229 -100
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 29 -188 229 -172
rect 287 -138 487 -100
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 287 -188 487 -172
rect 545 -138 745 -100
rect 545 -172 561 -138
rect 729 -172 745 -138
rect 545 -188 745 -172
rect 803 -138 1003 -100
rect 803 -172 819 -138
rect 987 -172 1003 -138
rect 803 -188 1003 -172
rect 1061 -138 1261 -100
rect 1061 -172 1077 -138
rect 1245 -172 1261 -138
rect 1061 -188 1261 -172
rect 1319 -138 1519 -100
rect 1319 -172 1335 -138
rect 1503 -172 1519 -138
rect 1319 -188 1519 -172
rect 1577 -138 1777 -100
rect 1577 -172 1593 -138
rect 1761 -172 1777 -138
rect 1577 -188 1777 -172
rect 1835 -138 2035 -100
rect 1835 -172 1851 -138
rect 2019 -172 2035 -138
rect 1835 -188 2035 -172
rect 2093 -138 2293 -100
rect 2093 -172 2109 -138
rect 2277 -172 2293 -138
rect 2093 -188 2293 -172
rect 2351 -138 2551 -100
rect 2351 -172 2367 -138
rect 2535 -172 2551 -138
rect 2351 -188 2551 -172
<< polycont >>
rect -2535 138 -2367 172
rect -2277 138 -2109 172
rect -2019 138 -1851 172
rect -1761 138 -1593 172
rect -1503 138 -1335 172
rect -1245 138 -1077 172
rect -987 138 -819 172
rect -729 138 -561 172
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect 561 138 729 172
rect 819 138 987 172
rect 1077 138 1245 172
rect 1335 138 1503 172
rect 1593 138 1761 172
rect 1851 138 2019 172
rect 2109 138 2277 172
rect 2367 138 2535 172
rect -2535 -172 -2367 -138
rect -2277 -172 -2109 -138
rect -2019 -172 -1851 -138
rect -1761 -172 -1593 -138
rect -1503 -172 -1335 -138
rect -1245 -172 -1077 -138
rect -987 -172 -819 -138
rect -729 -172 -561 -138
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
rect 561 -172 729 -138
rect 819 -172 987 -138
rect 1077 -172 1245 -138
rect 1335 -172 1503 -138
rect 1593 -172 1761 -138
rect 1851 -172 2019 -138
rect 2109 -172 2277 -138
rect 2367 -172 2535 -138
<< locali >>
rect -2711 240 -2615 274
rect 2615 240 2711 274
rect 2677 178 2711 240
rect -2551 138 -2535 172
rect -2367 138 -2351 172
rect -2293 138 -2277 172
rect -2109 138 -2093 172
rect -2035 138 -2019 172
rect -1851 138 -1835 172
rect -1777 138 -1761 172
rect -1593 138 -1577 172
rect -1519 138 -1503 172
rect -1335 138 -1319 172
rect -1261 138 -1245 172
rect -1077 138 -1061 172
rect -1003 138 -987 172
rect -819 138 -803 172
rect -745 138 -729 172
rect -561 138 -545 172
rect -487 138 -471 172
rect -303 138 -287 172
rect -229 138 -213 172
rect -45 138 -29 172
rect 29 138 45 172
rect 213 138 229 172
rect 287 138 303 172
rect 471 138 487 172
rect 545 138 561 172
rect 729 138 745 172
rect 803 138 819 172
rect 987 138 1003 172
rect 1061 138 1077 172
rect 1245 138 1261 172
rect 1319 138 1335 172
rect 1503 138 1519 172
rect 1577 138 1593 172
rect 1761 138 1777 172
rect 1835 138 1851 172
rect 2019 138 2035 172
rect 2093 138 2109 172
rect 2277 138 2293 172
rect 2351 138 2367 172
rect 2535 138 2551 172
rect -2597 88 -2563 104
rect -2597 -104 -2563 -88
rect -2339 88 -2305 104
rect -2339 -104 -2305 -88
rect -2081 88 -2047 104
rect -2081 -104 -2047 -88
rect -1823 88 -1789 104
rect -1823 -104 -1789 -88
rect -1565 88 -1531 104
rect -1565 -104 -1531 -88
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect 1531 88 1565 104
rect 1531 -104 1565 -88
rect 1789 88 1823 104
rect 1789 -104 1823 -88
rect 2047 88 2081 104
rect 2047 -104 2081 -88
rect 2305 88 2339 104
rect 2305 -104 2339 -88
rect 2563 88 2597 104
rect 2563 -104 2597 -88
rect -2551 -172 -2535 -138
rect -2367 -172 -2351 -138
rect -2293 -172 -2277 -138
rect -2109 -172 -2093 -138
rect -2035 -172 -2019 -138
rect -1851 -172 -1835 -138
rect -1777 -172 -1761 -138
rect -1593 -172 -1577 -138
rect -1519 -172 -1503 -138
rect -1335 -172 -1319 -138
rect -1261 -172 -1245 -138
rect -1077 -172 -1061 -138
rect -1003 -172 -987 -138
rect -819 -172 -803 -138
rect -745 -172 -729 -138
rect -561 -172 -545 -138
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 545 -172 561 -138
rect 729 -172 745 -138
rect 803 -172 819 -138
rect 987 -172 1003 -138
rect 1061 -172 1077 -138
rect 1245 -172 1261 -138
rect 1319 -172 1335 -138
rect 1503 -172 1519 -138
rect 1577 -172 1593 -138
rect 1761 -172 1777 -138
rect 1835 -172 1851 -138
rect 2019 -172 2035 -138
rect 2093 -172 2109 -138
rect 2277 -172 2293 -138
rect 2351 -172 2367 -138
rect 2535 -172 2551 -138
rect 2677 -240 2711 -178
rect -2711 -274 -2615 -240
rect 2615 -274 2711 -240
<< viali >>
rect -2711 178 -2677 240
rect -2711 -178 -2677 178
rect -2510 138 -2392 172
rect -2252 138 -2134 172
rect -1994 138 -1876 172
rect -1736 138 -1618 172
rect -1478 138 -1360 172
rect -1220 138 -1102 172
rect -962 138 -844 172
rect -704 138 -586 172
rect -446 138 -328 172
rect -188 138 -70 172
rect 70 138 188 172
rect 328 138 446 172
rect 586 138 704 172
rect 844 138 962 172
rect 1102 138 1220 172
rect 1360 138 1478 172
rect 1618 138 1736 172
rect 1876 138 1994 172
rect 2134 138 2252 172
rect 2392 138 2510 172
rect -2597 -88 -2563 88
rect -2339 -88 -2305 88
rect -2081 -88 -2047 88
rect -1823 -88 -1789 88
rect -1565 -88 -1531 88
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect 1531 -88 1565 88
rect 1789 -88 1823 88
rect 2047 -88 2081 88
rect 2305 -88 2339 88
rect 2563 -88 2597 88
rect -2510 -172 -2392 -138
rect -2252 -172 -2134 -138
rect -1994 -172 -1876 -138
rect -1736 -172 -1618 -138
rect -1478 -172 -1360 -138
rect -1220 -172 -1102 -138
rect -962 -172 -844 -138
rect -704 -172 -586 -138
rect -446 -172 -328 -138
rect -188 -172 -70 -138
rect 70 -172 188 -138
rect 328 -172 446 -138
rect 586 -172 704 -138
rect 844 -172 962 -138
rect 1102 -172 1220 -138
rect 1360 -172 1478 -138
rect 1618 -172 1736 -138
rect 1876 -172 1994 -138
rect 2134 -172 2252 -138
rect 2392 -172 2510 -138
rect -2711 -240 -2677 -178
<< metal1 >>
rect -2717 240 -2671 252
rect -2717 -240 -2711 240
rect -2677 -240 -2671 240
rect -2522 172 -2380 178
rect -2522 138 -2510 172
rect -2392 138 -2380 172
rect -2522 132 -2380 138
rect -2264 172 -2122 178
rect -2264 138 -2252 172
rect -2134 138 -2122 172
rect -2264 132 -2122 138
rect -2006 172 -1864 178
rect -2006 138 -1994 172
rect -1876 138 -1864 172
rect -2006 132 -1864 138
rect -1748 172 -1606 178
rect -1748 138 -1736 172
rect -1618 138 -1606 172
rect -1748 132 -1606 138
rect -1490 172 -1348 178
rect -1490 138 -1478 172
rect -1360 138 -1348 172
rect -1490 132 -1348 138
rect -1232 172 -1090 178
rect -1232 138 -1220 172
rect -1102 138 -1090 172
rect -1232 132 -1090 138
rect -974 172 -832 178
rect -974 138 -962 172
rect -844 138 -832 172
rect -974 132 -832 138
rect -716 172 -574 178
rect -716 138 -704 172
rect -586 138 -574 172
rect -716 132 -574 138
rect -458 172 -316 178
rect -458 138 -446 172
rect -328 138 -316 172
rect -458 132 -316 138
rect -200 172 -58 178
rect -200 138 -188 172
rect -70 138 -58 172
rect -200 132 -58 138
rect 58 172 200 178
rect 58 138 70 172
rect 188 138 200 172
rect 58 132 200 138
rect 316 172 458 178
rect 316 138 328 172
rect 446 138 458 172
rect 316 132 458 138
rect 574 172 716 178
rect 574 138 586 172
rect 704 138 716 172
rect 574 132 716 138
rect 832 172 974 178
rect 832 138 844 172
rect 962 138 974 172
rect 832 132 974 138
rect 1090 172 1232 178
rect 1090 138 1102 172
rect 1220 138 1232 172
rect 1090 132 1232 138
rect 1348 172 1490 178
rect 1348 138 1360 172
rect 1478 138 1490 172
rect 1348 132 1490 138
rect 1606 172 1748 178
rect 1606 138 1618 172
rect 1736 138 1748 172
rect 1606 132 1748 138
rect 1864 172 2006 178
rect 1864 138 1876 172
rect 1994 138 2006 172
rect 1864 132 2006 138
rect 2122 172 2264 178
rect 2122 138 2134 172
rect 2252 138 2264 172
rect 2122 132 2264 138
rect 2380 172 2522 178
rect 2380 138 2392 172
rect 2510 138 2522 172
rect 2380 132 2522 138
rect -2603 88 -2557 100
rect -2603 -88 -2597 88
rect -2563 -88 -2557 88
rect -2603 -100 -2557 -88
rect -2345 88 -2299 100
rect -2345 -88 -2339 88
rect -2305 -88 -2299 88
rect -2345 -100 -2299 -88
rect -2087 88 -2041 100
rect -2087 -88 -2081 88
rect -2047 -88 -2041 88
rect -2087 -100 -2041 -88
rect -1829 88 -1783 100
rect -1829 -88 -1823 88
rect -1789 -88 -1783 88
rect -1829 -100 -1783 -88
rect -1571 88 -1525 100
rect -1571 -88 -1565 88
rect -1531 -88 -1525 88
rect -1571 -100 -1525 -88
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect 1525 88 1571 100
rect 1525 -88 1531 88
rect 1565 -88 1571 88
rect 1525 -100 1571 -88
rect 1783 88 1829 100
rect 1783 -88 1789 88
rect 1823 -88 1829 88
rect 1783 -100 1829 -88
rect 2041 88 2087 100
rect 2041 -88 2047 88
rect 2081 -88 2087 88
rect 2041 -100 2087 -88
rect 2299 88 2345 100
rect 2299 -88 2305 88
rect 2339 -88 2345 88
rect 2299 -100 2345 -88
rect 2557 88 2603 100
rect 2557 -88 2563 88
rect 2597 -88 2603 88
rect 2557 -100 2603 -88
rect -2522 -138 -2380 -132
rect -2522 -172 -2510 -138
rect -2392 -172 -2380 -138
rect -2522 -178 -2380 -172
rect -2264 -138 -2122 -132
rect -2264 -172 -2252 -138
rect -2134 -172 -2122 -138
rect -2264 -178 -2122 -172
rect -2006 -138 -1864 -132
rect -2006 -172 -1994 -138
rect -1876 -172 -1864 -138
rect -2006 -178 -1864 -172
rect -1748 -138 -1606 -132
rect -1748 -172 -1736 -138
rect -1618 -172 -1606 -138
rect -1748 -178 -1606 -172
rect -1490 -138 -1348 -132
rect -1490 -172 -1478 -138
rect -1360 -172 -1348 -138
rect -1490 -178 -1348 -172
rect -1232 -138 -1090 -132
rect -1232 -172 -1220 -138
rect -1102 -172 -1090 -138
rect -1232 -178 -1090 -172
rect -974 -138 -832 -132
rect -974 -172 -962 -138
rect -844 -172 -832 -138
rect -974 -178 -832 -172
rect -716 -138 -574 -132
rect -716 -172 -704 -138
rect -586 -172 -574 -138
rect -716 -178 -574 -172
rect -458 -138 -316 -132
rect -458 -172 -446 -138
rect -328 -172 -316 -138
rect -458 -178 -316 -172
rect -200 -138 -58 -132
rect -200 -172 -188 -138
rect -70 -172 -58 -138
rect -200 -178 -58 -172
rect 58 -138 200 -132
rect 58 -172 70 -138
rect 188 -172 200 -138
rect 58 -178 200 -172
rect 316 -138 458 -132
rect 316 -172 328 -138
rect 446 -172 458 -138
rect 316 -178 458 -172
rect 574 -138 716 -132
rect 574 -172 586 -138
rect 704 -172 716 -138
rect 574 -178 716 -172
rect 832 -138 974 -132
rect 832 -172 844 -138
rect 962 -172 974 -138
rect 832 -178 974 -172
rect 1090 -138 1232 -132
rect 1090 -172 1102 -138
rect 1220 -172 1232 -138
rect 1090 -178 1232 -172
rect 1348 -138 1490 -132
rect 1348 -172 1360 -138
rect 1478 -172 1490 -138
rect 1348 -178 1490 -172
rect 1606 -138 1748 -132
rect 1606 -172 1618 -138
rect 1736 -172 1748 -138
rect 1606 -178 1748 -172
rect 1864 -138 2006 -132
rect 1864 -172 1876 -138
rect 1994 -172 2006 -138
rect 1864 -178 2006 -172
rect 2122 -138 2264 -132
rect 2122 -172 2134 -138
rect 2252 -172 2264 -138
rect 2122 -178 2264 -172
rect 2380 -138 2522 -132
rect 2380 -172 2392 -138
rect 2510 -172 2522 -138
rect 2380 -178 2522 -172
rect -2717 -252 -2671 -240
<< properties >>
string FIXED_BBOX -2694 -257 2694 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 100 viagt 0
<< end >>
