magic
tech sky130A
magscale 1 2
timestamp 1675896495
<< metal4 >>
rect -2869 67839 2869 67880
rect -2869 62721 2613 67839
rect 2849 62721 2869 67839
rect -2869 62680 2869 62721
rect -2869 62399 2869 62440
rect -2869 57281 2613 62399
rect 2849 57281 2869 62399
rect -2869 57240 2869 57281
rect -2869 56959 2869 57000
rect -2869 51841 2613 56959
rect 2849 51841 2869 56959
rect -2869 51800 2869 51841
rect -2869 51519 2869 51560
rect -2869 46401 2613 51519
rect 2849 46401 2869 51519
rect -2869 46360 2869 46401
rect -2869 46079 2869 46120
rect -2869 40961 2613 46079
rect 2849 40961 2869 46079
rect -2869 40920 2869 40961
rect -2869 40639 2869 40680
rect -2869 35521 2613 40639
rect 2849 35521 2869 40639
rect -2869 35480 2869 35521
rect -2869 35199 2869 35240
rect -2869 30081 2613 35199
rect 2849 30081 2869 35199
rect -2869 30040 2869 30081
rect -2869 29759 2869 29800
rect -2869 24641 2613 29759
rect 2849 24641 2869 29759
rect -2869 24600 2869 24641
rect -2869 24319 2869 24360
rect -2869 19201 2613 24319
rect 2849 19201 2869 24319
rect -2869 19160 2869 19201
rect -2869 18879 2869 18920
rect -2869 13761 2613 18879
rect 2849 13761 2869 18879
rect -2869 13720 2869 13761
rect -2869 13439 2869 13480
rect -2869 8321 2613 13439
rect 2849 8321 2869 13439
rect -2869 8280 2869 8321
rect -2869 7999 2869 8040
rect -2869 2881 2613 7999
rect 2849 2881 2869 7999
rect -2869 2840 2869 2881
rect -2869 2559 2869 2600
rect -2869 -2559 2613 2559
rect 2849 -2559 2869 2559
rect -2869 -2600 2869 -2559
rect -2869 -2881 2869 -2840
rect -2869 -7999 2613 -2881
rect 2849 -7999 2869 -2881
rect -2869 -8040 2869 -7999
rect -2869 -8321 2869 -8280
rect -2869 -13439 2613 -8321
rect 2849 -13439 2869 -8321
rect -2869 -13480 2869 -13439
rect -2869 -13761 2869 -13720
rect -2869 -18879 2613 -13761
rect 2849 -18879 2869 -13761
rect -2869 -18920 2869 -18879
rect -2869 -19201 2869 -19160
rect -2869 -24319 2613 -19201
rect 2849 -24319 2869 -19201
rect -2869 -24360 2869 -24319
rect -2869 -24641 2869 -24600
rect -2869 -29759 2613 -24641
rect 2849 -29759 2869 -24641
rect -2869 -29800 2869 -29759
rect -2869 -30081 2869 -30040
rect -2869 -35199 2613 -30081
rect 2849 -35199 2869 -30081
rect -2869 -35240 2869 -35199
rect -2869 -35521 2869 -35480
rect -2869 -40639 2613 -35521
rect 2849 -40639 2869 -35521
rect -2869 -40680 2869 -40639
rect -2869 -40961 2869 -40920
rect -2869 -46079 2613 -40961
rect 2849 -46079 2869 -40961
rect -2869 -46120 2869 -46079
rect -2869 -46401 2869 -46360
rect -2869 -51519 2613 -46401
rect 2849 -51519 2869 -46401
rect -2869 -51560 2869 -51519
rect -2869 -51841 2869 -51800
rect -2869 -56959 2613 -51841
rect 2849 -56959 2869 -51841
rect -2869 -57000 2869 -56959
rect -2869 -57281 2869 -57240
rect -2869 -62399 2613 -57281
rect 2849 -62399 2869 -57281
rect -2869 -62440 2869 -62399
rect -2869 -62721 2869 -62680
rect -2869 -67839 2613 -62721
rect 2849 -67839 2869 -62721
rect -2869 -67880 2869 -67839
<< via4 >>
rect 2613 62721 2849 67839
rect 2613 57281 2849 62399
rect 2613 51841 2849 56959
rect 2613 46401 2849 51519
rect 2613 40961 2849 46079
rect 2613 35521 2849 40639
rect 2613 30081 2849 35199
rect 2613 24641 2849 29759
rect 2613 19201 2849 24319
rect 2613 13761 2849 18879
rect 2613 8321 2849 13439
rect 2613 2881 2849 7999
rect 2613 -2559 2849 2559
rect 2613 -7999 2849 -2881
rect 2613 -13439 2849 -8321
rect 2613 -18879 2849 -13761
rect 2613 -24319 2849 -19201
rect 2613 -29759 2849 -24641
rect 2613 -35199 2849 -30081
rect 2613 -40639 2849 -35521
rect 2613 -46079 2849 -40961
rect 2613 -51519 2849 -46401
rect 2613 -56959 2849 -51841
rect 2613 -62399 2849 -57281
rect 2613 -67839 2849 -62721
<< mimcap2 >>
rect -2789 67760 2251 67800
rect -2789 62800 -2749 67760
rect 2211 62800 2251 67760
rect -2789 62760 2251 62800
rect -2789 62320 2251 62360
rect -2789 57360 -2749 62320
rect 2211 57360 2251 62320
rect -2789 57320 2251 57360
rect -2789 56880 2251 56920
rect -2789 51920 -2749 56880
rect 2211 51920 2251 56880
rect -2789 51880 2251 51920
rect -2789 51440 2251 51480
rect -2789 46480 -2749 51440
rect 2211 46480 2251 51440
rect -2789 46440 2251 46480
rect -2789 46000 2251 46040
rect -2789 41040 -2749 46000
rect 2211 41040 2251 46000
rect -2789 41000 2251 41040
rect -2789 40560 2251 40600
rect -2789 35600 -2749 40560
rect 2211 35600 2251 40560
rect -2789 35560 2251 35600
rect -2789 35120 2251 35160
rect -2789 30160 -2749 35120
rect 2211 30160 2251 35120
rect -2789 30120 2251 30160
rect -2789 29680 2251 29720
rect -2789 24720 -2749 29680
rect 2211 24720 2251 29680
rect -2789 24680 2251 24720
rect -2789 24240 2251 24280
rect -2789 19280 -2749 24240
rect 2211 19280 2251 24240
rect -2789 19240 2251 19280
rect -2789 18800 2251 18840
rect -2789 13840 -2749 18800
rect 2211 13840 2251 18800
rect -2789 13800 2251 13840
rect -2789 13360 2251 13400
rect -2789 8400 -2749 13360
rect 2211 8400 2251 13360
rect -2789 8360 2251 8400
rect -2789 7920 2251 7960
rect -2789 2960 -2749 7920
rect 2211 2960 2251 7920
rect -2789 2920 2251 2960
rect -2789 2480 2251 2520
rect -2789 -2480 -2749 2480
rect 2211 -2480 2251 2480
rect -2789 -2520 2251 -2480
rect -2789 -2960 2251 -2920
rect -2789 -7920 -2749 -2960
rect 2211 -7920 2251 -2960
rect -2789 -7960 2251 -7920
rect -2789 -8400 2251 -8360
rect -2789 -13360 -2749 -8400
rect 2211 -13360 2251 -8400
rect -2789 -13400 2251 -13360
rect -2789 -13840 2251 -13800
rect -2789 -18800 -2749 -13840
rect 2211 -18800 2251 -13840
rect -2789 -18840 2251 -18800
rect -2789 -19280 2251 -19240
rect -2789 -24240 -2749 -19280
rect 2211 -24240 2251 -19280
rect -2789 -24280 2251 -24240
rect -2789 -24720 2251 -24680
rect -2789 -29680 -2749 -24720
rect 2211 -29680 2251 -24720
rect -2789 -29720 2251 -29680
rect -2789 -30160 2251 -30120
rect -2789 -35120 -2749 -30160
rect 2211 -35120 2251 -30160
rect -2789 -35160 2251 -35120
rect -2789 -35600 2251 -35560
rect -2789 -40560 -2749 -35600
rect 2211 -40560 2251 -35600
rect -2789 -40600 2251 -40560
rect -2789 -41040 2251 -41000
rect -2789 -46000 -2749 -41040
rect 2211 -46000 2251 -41040
rect -2789 -46040 2251 -46000
rect -2789 -46480 2251 -46440
rect -2789 -51440 -2749 -46480
rect 2211 -51440 2251 -46480
rect -2789 -51480 2251 -51440
rect -2789 -51920 2251 -51880
rect -2789 -56880 -2749 -51920
rect 2211 -56880 2251 -51920
rect -2789 -56920 2251 -56880
rect -2789 -57360 2251 -57320
rect -2789 -62320 -2749 -57360
rect 2211 -62320 2251 -57360
rect -2789 -62360 2251 -62320
rect -2789 -62800 2251 -62760
rect -2789 -67760 -2749 -62800
rect 2211 -67760 2251 -62800
rect -2789 -67800 2251 -67760
<< mimcap2contact >>
rect -2749 62800 2211 67760
rect -2749 57360 2211 62320
rect -2749 51920 2211 56880
rect -2749 46480 2211 51440
rect -2749 41040 2211 46000
rect -2749 35600 2211 40560
rect -2749 30160 2211 35120
rect -2749 24720 2211 29680
rect -2749 19280 2211 24240
rect -2749 13840 2211 18800
rect -2749 8400 2211 13360
rect -2749 2960 2211 7920
rect -2749 -2480 2211 2480
rect -2749 -7920 2211 -2960
rect -2749 -13360 2211 -8400
rect -2749 -18800 2211 -13840
rect -2749 -24240 2211 -19280
rect -2749 -29680 2211 -24720
rect -2749 -35120 2211 -30160
rect -2749 -40560 2211 -35600
rect -2749 -46000 2211 -41040
rect -2749 -51440 2211 -46480
rect -2749 -56880 2211 -51920
rect -2749 -62320 2211 -57360
rect -2749 -67760 2211 -62800
<< metal5 >>
rect -429 67784 -109 68000
rect 2571 67839 2891 68000
rect -2773 67760 2235 67784
rect -2773 62800 -2749 67760
rect 2211 62800 2235 67760
rect -2773 62776 2235 62800
rect -429 62344 -109 62776
rect 2571 62721 2613 67839
rect 2849 62721 2891 67839
rect 2571 62399 2891 62721
rect -2773 62320 2235 62344
rect -2773 57360 -2749 62320
rect 2211 57360 2235 62320
rect -2773 57336 2235 57360
rect -429 56904 -109 57336
rect 2571 57281 2613 62399
rect 2849 57281 2891 62399
rect 2571 56959 2891 57281
rect -2773 56880 2235 56904
rect -2773 51920 -2749 56880
rect 2211 51920 2235 56880
rect -2773 51896 2235 51920
rect -429 51464 -109 51896
rect 2571 51841 2613 56959
rect 2849 51841 2891 56959
rect 2571 51519 2891 51841
rect -2773 51440 2235 51464
rect -2773 46480 -2749 51440
rect 2211 46480 2235 51440
rect -2773 46456 2235 46480
rect -429 46024 -109 46456
rect 2571 46401 2613 51519
rect 2849 46401 2891 51519
rect 2571 46079 2891 46401
rect -2773 46000 2235 46024
rect -2773 41040 -2749 46000
rect 2211 41040 2235 46000
rect -2773 41016 2235 41040
rect -429 40584 -109 41016
rect 2571 40961 2613 46079
rect 2849 40961 2891 46079
rect 2571 40639 2891 40961
rect -2773 40560 2235 40584
rect -2773 35600 -2749 40560
rect 2211 35600 2235 40560
rect -2773 35576 2235 35600
rect -429 35144 -109 35576
rect 2571 35521 2613 40639
rect 2849 35521 2891 40639
rect 2571 35199 2891 35521
rect -2773 35120 2235 35144
rect -2773 30160 -2749 35120
rect 2211 30160 2235 35120
rect -2773 30136 2235 30160
rect -429 29704 -109 30136
rect 2571 30081 2613 35199
rect 2849 30081 2891 35199
rect 2571 29759 2891 30081
rect -2773 29680 2235 29704
rect -2773 24720 -2749 29680
rect 2211 24720 2235 29680
rect -2773 24696 2235 24720
rect -429 24264 -109 24696
rect 2571 24641 2613 29759
rect 2849 24641 2891 29759
rect 2571 24319 2891 24641
rect -2773 24240 2235 24264
rect -2773 19280 -2749 24240
rect 2211 19280 2235 24240
rect -2773 19256 2235 19280
rect -429 18824 -109 19256
rect 2571 19201 2613 24319
rect 2849 19201 2891 24319
rect 2571 18879 2891 19201
rect -2773 18800 2235 18824
rect -2773 13840 -2749 18800
rect 2211 13840 2235 18800
rect -2773 13816 2235 13840
rect -429 13384 -109 13816
rect 2571 13761 2613 18879
rect 2849 13761 2891 18879
rect 2571 13439 2891 13761
rect -2773 13360 2235 13384
rect -2773 8400 -2749 13360
rect 2211 8400 2235 13360
rect -2773 8376 2235 8400
rect -429 7944 -109 8376
rect 2571 8321 2613 13439
rect 2849 8321 2891 13439
rect 2571 7999 2891 8321
rect -2773 7920 2235 7944
rect -2773 2960 -2749 7920
rect 2211 2960 2235 7920
rect -2773 2936 2235 2960
rect -429 2504 -109 2936
rect 2571 2881 2613 7999
rect 2849 2881 2891 7999
rect 2571 2559 2891 2881
rect -2773 2480 2235 2504
rect -2773 -2480 -2749 2480
rect 2211 -2480 2235 2480
rect -2773 -2504 2235 -2480
rect -429 -2936 -109 -2504
rect 2571 -2559 2613 2559
rect 2849 -2559 2891 2559
rect 2571 -2881 2891 -2559
rect -2773 -2960 2235 -2936
rect -2773 -7920 -2749 -2960
rect 2211 -7920 2235 -2960
rect -2773 -7944 2235 -7920
rect -429 -8376 -109 -7944
rect 2571 -7999 2613 -2881
rect 2849 -7999 2891 -2881
rect 2571 -8321 2891 -7999
rect -2773 -8400 2235 -8376
rect -2773 -13360 -2749 -8400
rect 2211 -13360 2235 -8400
rect -2773 -13384 2235 -13360
rect -429 -13816 -109 -13384
rect 2571 -13439 2613 -8321
rect 2849 -13439 2891 -8321
rect 2571 -13761 2891 -13439
rect -2773 -13840 2235 -13816
rect -2773 -18800 -2749 -13840
rect 2211 -18800 2235 -13840
rect -2773 -18824 2235 -18800
rect -429 -19256 -109 -18824
rect 2571 -18879 2613 -13761
rect 2849 -18879 2891 -13761
rect 2571 -19201 2891 -18879
rect -2773 -19280 2235 -19256
rect -2773 -24240 -2749 -19280
rect 2211 -24240 2235 -19280
rect -2773 -24264 2235 -24240
rect -429 -24696 -109 -24264
rect 2571 -24319 2613 -19201
rect 2849 -24319 2891 -19201
rect 2571 -24641 2891 -24319
rect -2773 -24720 2235 -24696
rect -2773 -29680 -2749 -24720
rect 2211 -29680 2235 -24720
rect -2773 -29704 2235 -29680
rect -429 -30136 -109 -29704
rect 2571 -29759 2613 -24641
rect 2849 -29759 2891 -24641
rect 2571 -30081 2891 -29759
rect -2773 -30160 2235 -30136
rect -2773 -35120 -2749 -30160
rect 2211 -35120 2235 -30160
rect -2773 -35144 2235 -35120
rect -429 -35576 -109 -35144
rect 2571 -35199 2613 -30081
rect 2849 -35199 2891 -30081
rect 2571 -35521 2891 -35199
rect -2773 -35600 2235 -35576
rect -2773 -40560 -2749 -35600
rect 2211 -40560 2235 -35600
rect -2773 -40584 2235 -40560
rect -429 -41016 -109 -40584
rect 2571 -40639 2613 -35521
rect 2849 -40639 2891 -35521
rect 2571 -40961 2891 -40639
rect -2773 -41040 2235 -41016
rect -2773 -46000 -2749 -41040
rect 2211 -46000 2235 -41040
rect -2773 -46024 2235 -46000
rect -429 -46456 -109 -46024
rect 2571 -46079 2613 -40961
rect 2849 -46079 2891 -40961
rect 2571 -46401 2891 -46079
rect -2773 -46480 2235 -46456
rect -2773 -51440 -2749 -46480
rect 2211 -51440 2235 -46480
rect -2773 -51464 2235 -51440
rect -429 -51896 -109 -51464
rect 2571 -51519 2613 -46401
rect 2849 -51519 2891 -46401
rect 2571 -51841 2891 -51519
rect -2773 -51920 2235 -51896
rect -2773 -56880 -2749 -51920
rect 2211 -56880 2235 -51920
rect -2773 -56904 2235 -56880
rect -429 -57336 -109 -56904
rect 2571 -56959 2613 -51841
rect 2849 -56959 2891 -51841
rect 2571 -57281 2891 -56959
rect -2773 -57360 2235 -57336
rect -2773 -62320 -2749 -57360
rect 2211 -62320 2235 -57360
rect -2773 -62344 2235 -62320
rect -429 -62776 -109 -62344
rect 2571 -62399 2613 -57281
rect 2849 -62399 2891 -57281
rect 2571 -62721 2891 -62399
rect -2773 -62800 2235 -62776
rect -2773 -67760 -2749 -62800
rect 2211 -67760 2235 -62800
rect -2773 -67784 2235 -67760
rect -429 -68000 -109 -67784
rect 2571 -67839 2613 -62721
rect 2849 -67839 2891 -62721
rect 2571 -68000 2891 -67839
<< properties >>
string FIXED_BBOX -2869 62680 2331 67880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.2 l 25.2 val 1.289k carea 2.00 cperi 0.19 nx 1 ny 25 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
