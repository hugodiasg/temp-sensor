** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator_tb-tran.sch
**.subckt ask-modulator_tb-tran
Vdd vd GND 3.3
Vin in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 100ns 200ns)
x1 vd out in GND ask-modulator
**** begin user architecture code


*.tran 0.3n 110n
*.tran 0.5n 200n
.tran 1n 1000n
.control
destroy all
run
let id =-i(vdd)
let z_rlc= (vd-out)/id
let z_nmos=out/id
let z_out=z_rlc*z_nmos/(z_rlc+z_nmos)
plot z_out
plot id
plot in
plot out
let S=abs(id*(vd-out))+abs(id*out)
plot s
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  ask-modulator.sym # of pins=4
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sch
.subckt ask-modulator  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XM2 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=24 L=24 MF=3 m=3
XR0 out vd gnd sky130_fd_pr__res_high_po_5p73 L=0.56 mult=4 m=4
x1 vd out l0
**** begin user architecture code

*X0 out.t4 out.t5 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X1 out in.t0 gnd gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p
*+ ps=1.798e+07u w=0u l=0u
*X2 out.t0 out.t1 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X3 out.t2 out.t3 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 out.n2 out 3.44
R1 out.n3 out 2.874
R2 out out.n2 1.395
R3 out.n0 out.t5 0.485
R4 out.n1 out.n0 0.484
R5 out.n3 out.t0 0.146
R6 out.n2 out.n1 0.122
R7 out.t2 out.t4 0.064
R8 out.t0 out.t2 0.064
R9 out out.n3 0.042
R10 out.n0 out.t3 0.023
R11 out.n1 out.t1 0.001
R12 in in.t0 446.69
C0 in gnd 0.98fF
C1 out in 0.05fF
C2 out gnd 3.40fF
C3 out.t3 0 8.30fF
C4 out.t5 0 11.92fF
C5 out.n0 0 4.15fF $ **FLOATING
C6 out.t1 0 5.68fF
C7 out.n1 0 6.72fF $ **FLOATING
C8 out.n2 0 20.76fF $ **FLOATING
C9 out.t4 0 18.71fF
C10 out.t2 0 18.76fF
C11 out.t0 0 19.44fF
C12 out.n3 0 15.11fF $ **FLOATING
C13 out 0 314.11fF
C14 gnd 0 12.33fF
C15 in 0 1.73fF

**** end user architecture code
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym # of
*+ pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sch
.subckt l0  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.006n m=1
Cs1 p1 net1 10.86f m=1
Cs2 p2 net2 11.96f m=1
Rs1 net1 GND 114.5 m=1
Rs2 net2 GND -66.9 m=1
R1 p2 net3 5.426 m=1
.ends

.GLOBAL GND
.end
