magic
tech sky130A
magscale 1 2
timestamp 1643669011
<< pwell >>
rect -844 -678 844 678
<< mvnmos >>
rect -616 -420 -416 420
rect -358 -420 -158 420
rect -100 -420 100 420
rect 158 -420 358 420
rect 416 -420 616 420
<< mvndiff >>
rect -674 408 -616 420
rect -674 -408 -662 408
rect -628 -408 -616 408
rect -674 -420 -616 -408
rect -416 408 -358 420
rect -416 -408 -404 408
rect -370 -408 -358 408
rect -416 -420 -358 -408
rect -158 408 -100 420
rect -158 -408 -146 408
rect -112 -408 -100 408
rect -158 -420 -100 -408
rect 100 408 158 420
rect 100 -408 112 408
rect 146 -408 158 408
rect 100 -420 158 -408
rect 358 408 416 420
rect 358 -408 370 408
rect 404 -408 416 408
rect 358 -420 416 -408
rect 616 408 674 420
rect 616 -408 628 408
rect 662 -408 674 408
rect 616 -420 674 -408
<< mvndiffc >>
rect -662 -408 -628 408
rect -404 -408 -370 408
rect -146 -408 -112 408
rect 112 -408 146 408
rect 370 -408 404 408
rect 628 -408 662 408
<< mvpsubdiff >>
rect -808 630 808 642
rect -808 596 -700 630
rect 700 596 808 630
rect -808 584 808 596
rect -808 534 -750 584
rect -808 -534 -796 534
rect -762 -534 -750 534
rect 750 534 808 584
rect -808 -584 -750 -534
rect 750 -534 762 534
rect 796 -534 808 534
rect 750 -584 808 -534
rect -808 -596 808 -584
rect -808 -630 -700 -596
rect 700 -630 808 -596
rect -808 -642 808 -630
<< mvpsubdiffcont >>
rect -700 596 700 630
rect -796 -534 -762 534
rect 762 -534 796 534
rect -700 -630 700 -596
<< poly >>
rect -616 492 -416 508
rect -616 458 -600 492
rect -432 458 -416 492
rect -616 420 -416 458
rect -358 492 -158 508
rect -358 458 -342 492
rect -174 458 -158 492
rect -358 420 -158 458
rect -100 492 100 508
rect -100 458 -84 492
rect 84 458 100 492
rect -100 420 100 458
rect 158 492 358 508
rect 158 458 174 492
rect 342 458 358 492
rect 158 420 358 458
rect 416 492 616 508
rect 416 458 432 492
rect 600 458 616 492
rect 416 420 616 458
rect -616 -458 -416 -420
rect -616 -492 -600 -458
rect -432 -492 -416 -458
rect -616 -508 -416 -492
rect -358 -458 -158 -420
rect -358 -492 -342 -458
rect -174 -492 -158 -458
rect -358 -508 -158 -492
rect -100 -458 100 -420
rect -100 -492 -84 -458
rect 84 -492 100 -458
rect -100 -508 100 -492
rect 158 -458 358 -420
rect 158 -492 174 -458
rect 342 -492 358 -458
rect 158 -508 358 -492
rect 416 -458 616 -420
rect 416 -492 432 -458
rect 600 -492 616 -458
rect 416 -508 616 -492
<< polycont >>
rect -600 458 -432 492
rect -342 458 -174 492
rect -84 458 84 492
rect 174 458 342 492
rect 432 458 600 492
rect -600 -492 -432 -458
rect -342 -492 -174 -458
rect -84 -492 84 -458
rect 174 -492 342 -458
rect 432 -492 600 -458
<< locali >>
rect -796 596 -700 630
rect 700 596 796 630
rect -796 534 -762 596
rect 762 534 796 596
rect -616 458 -600 492
rect -432 458 -416 492
rect -358 458 -342 492
rect -174 458 -158 492
rect -100 458 -84 492
rect 84 458 100 492
rect 158 458 174 492
rect 342 458 358 492
rect 416 458 432 492
rect 600 458 616 492
rect -662 408 -628 424
rect -662 -424 -628 -408
rect -404 408 -370 424
rect -404 -424 -370 -408
rect -146 408 -112 424
rect -146 -424 -112 -408
rect 112 408 146 424
rect 112 -424 146 -408
rect 370 408 404 424
rect 370 -424 404 -408
rect 628 408 662 424
rect 628 -424 662 -408
rect -616 -492 -600 -458
rect -432 -492 -416 -458
rect -358 -492 -342 -458
rect -174 -492 -158 -458
rect -100 -492 -84 -458
rect 84 -492 100 -458
rect 158 -492 174 -458
rect 342 -492 358 -458
rect 416 -492 432 -458
rect 600 -492 616 -458
rect -796 -630 -762 -534
rect 762 -630 796 -534
<< viali >>
rect -600 458 -432 492
rect -342 458 -174 492
rect -84 458 84 492
rect 174 458 342 492
rect 432 458 600 492
rect -662 -17 -628 391
rect -404 -204 -370 204
rect -146 -17 -112 391
rect 112 -204 146 204
rect 370 -17 404 391
rect 628 -204 662 204
rect -600 -492 -432 -458
rect -342 -492 -174 -458
rect -84 -492 84 -458
rect 174 -492 342 -458
rect 432 -492 600 -458
rect -762 -630 -700 -596
rect -700 -630 700 -596
rect 700 -630 762 -596
<< metal1 >>
rect -612 492 -420 498
rect -612 458 -600 492
rect -432 458 -420 492
rect -612 452 -420 458
rect -354 492 -162 498
rect -354 458 -342 492
rect -174 458 -162 492
rect -354 452 -162 458
rect -96 492 96 498
rect -96 458 -84 492
rect 84 458 96 492
rect -96 452 96 458
rect 162 492 354 498
rect 162 458 174 492
rect 342 458 354 492
rect 162 452 354 458
rect 420 492 612 498
rect 420 458 432 492
rect 600 458 612 492
rect 420 452 612 458
rect -668 391 -622 403
rect -668 -17 -662 391
rect -628 -17 -622 391
rect -152 391 -106 403
rect -668 -29 -622 -17
rect -410 204 -364 216
rect -410 -204 -404 204
rect -370 -204 -364 204
rect -152 -17 -146 391
rect -112 -17 -106 391
rect 364 391 410 403
rect -152 -29 -106 -17
rect 106 204 152 216
rect -410 -216 -364 -204
rect 106 -204 112 204
rect 146 -204 152 204
rect 364 -17 370 391
rect 404 -17 410 391
rect 364 -29 410 -17
rect 622 204 668 216
rect 106 -216 152 -204
rect 622 -204 628 204
rect 662 -204 668 204
rect 622 -216 668 -204
rect -612 -458 -420 -452
rect -612 -492 -600 -458
rect -432 -492 -420 -458
rect -612 -498 -420 -492
rect -354 -458 -162 -452
rect -354 -492 -342 -458
rect -174 -492 -162 -458
rect -354 -498 -162 -492
rect -96 -458 96 -452
rect -96 -492 -84 -458
rect 84 -492 96 -458
rect -96 -498 96 -492
rect 162 -458 354 -452
rect 162 -492 174 -458
rect 342 -492 354 -458
rect 162 -498 354 -492
rect 420 -458 612 -452
rect 420 -492 432 -458
rect 600 -492 612 -458
rect 420 -498 612 -492
rect -774 -596 774 -590
rect -774 -630 -762 -596
rect 762 -630 774 -596
rect -774 -636 774 -630
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -779 -613 779 613
string parameters w 4.2 l 1.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 50 viadrn -50 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
