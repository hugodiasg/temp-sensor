magic
tech sky130A
timestamp 1700075225
<< pwell >>
rect -2098 -155 2098 155
<< nmos >>
rect -2000 -50 2000 50
<< ndiff >>
rect -2029 44 -2000 50
rect -2029 -44 -2023 44
rect -2006 -44 -2000 44
rect -2029 -50 -2000 -44
rect 2000 44 2029 50
rect 2000 -44 2006 44
rect 2023 -44 2029 44
rect 2000 -50 2029 -44
<< ndiffc >>
rect -2023 -44 -2006 44
rect 2006 -44 2023 44
<< psubdiff >>
rect -2080 120 -2032 137
rect 2032 120 2080 137
rect -2080 89 -2063 120
rect 2063 89 2080 120
rect -2080 -120 -2063 -89
rect 2063 -120 2080 -89
rect -2080 -137 -2032 -120
rect 2032 -137 2080 -120
<< psubdiffcont >>
rect -2032 120 2032 137
rect -2080 -89 -2063 89
rect 2063 -89 2080 89
rect -2032 -137 2032 -120
<< poly >>
rect -2000 86 2000 94
rect -2000 69 -1992 86
rect 1992 69 2000 86
rect -2000 50 2000 69
rect -2000 -69 2000 -50
rect -2000 -86 -1992 -69
rect 1992 -86 2000 -69
rect -2000 -94 2000 -86
<< polycont >>
rect -1992 69 1992 86
rect -1992 -86 1992 -69
<< locali >>
rect -2080 120 -2032 137
rect 2032 120 2080 137
rect -2080 89 -2063 120
rect 2063 89 2080 120
rect -2000 69 -1992 86
rect 1992 69 2000 86
rect -2023 44 -2006 52
rect -2023 -52 -2006 -44
rect 2006 44 2023 52
rect 2006 -52 2023 -44
rect -2000 -86 -1992 -69
rect 1992 -86 2000 -69
rect -2080 -120 -2063 -89
rect 2063 -120 2080 -89
rect -2080 -137 -2032 -120
rect 2032 -137 2080 -120
<< viali >>
rect -1992 69 1992 86
rect -2023 -44 -2006 44
rect 2006 -44 2023 44
rect -1992 -86 1992 -69
<< metal1 >>
rect -1998 86 1998 89
rect -1998 69 -1992 86
rect 1992 69 1998 86
rect -1998 66 1998 69
rect -2026 44 -2003 50
rect -2026 -44 -2023 44
rect -2006 -44 -2003 44
rect -2026 -50 -2003 -44
rect 2003 44 2026 50
rect 2003 -44 2006 44
rect 2023 -44 2026 44
rect 2003 -50 2026 -44
rect -1998 -69 1998 -66
rect -1998 -86 -1992 -69
rect 1992 -86 1998 -69
rect -1998 -89 1998 -86
<< properties >>
string FIXED_BBOX -2071 -128 2071 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 40 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
