magic
tech sky130A
magscale 1 2
timestamp 1657058092
<< nwell >>
rect 4340 2520 4932 3358
rect 4440 1400 5032 2238
rect 7640 850 7690 880
rect 7820 820 7846 1020
<< pmos >>
rect 4536 2739 4736 3139
rect 4636 1619 4836 2019
<< pdiff >>
rect 4478 3127 4536 3139
rect 4478 2751 4490 3127
rect 4524 2751 4536 3127
rect 4478 2739 4536 2751
rect 4736 3127 4794 3139
rect 4736 2751 4748 3127
rect 4782 2751 4794 3127
rect 4736 2739 4794 2751
rect 4578 2007 4636 2019
rect 4578 1631 4590 2007
rect 4624 1631 4636 2007
rect 4578 1619 4636 1631
rect 4836 2007 4894 2019
rect 4836 1631 4848 2007
rect 4882 1631 4894 2007
rect 4836 1619 4894 1631
<< pdiffc >>
rect 4490 2751 4524 3127
rect 4748 2751 4782 3127
rect 4590 1631 4624 2007
rect 4848 1631 4882 2007
<< psubdiff >>
rect 9086 130 9110 210
rect 9250 130 9274 210
<< nsubdiff >>
rect 4376 3288 4472 3322
rect 4800 3288 4896 3322
rect 4376 3226 4410 3288
rect 4862 3226 4896 3288
rect 4376 2590 4410 2652
rect 4862 2590 4896 2652
rect 4376 2556 4472 2590
rect 4800 2556 4896 2590
rect 4476 2168 4572 2202
rect 4900 2168 4996 2202
rect 4476 2106 4510 2168
rect 4962 2106 4996 2168
rect 4476 1470 4510 1532
rect 4962 1470 4996 1532
rect 4476 1436 4572 1470
rect 4900 1436 4996 1470
<< psubdiffcont >>
rect 9110 130 9250 210
<< nsubdiffcont >>
rect 4472 3288 4800 3322
rect 4376 2652 4410 3226
rect 4862 2652 4896 3226
rect 4472 2556 4800 2590
rect 4572 2168 4900 2202
rect 4476 1532 4510 2106
rect 4962 1532 4996 2106
rect 4572 1436 4900 1470
<< poly >>
rect 4536 3220 4736 3236
rect 4536 3186 4552 3220
rect 4720 3186 4736 3220
rect 4536 3139 4736 3186
rect 4536 2692 4736 2739
rect 4536 2658 4552 2692
rect 4720 2658 4736 2692
rect 4536 2642 4736 2658
rect 4636 2100 4836 2116
rect 4636 2066 4652 2100
rect 4820 2066 4836 2100
rect 4636 2019 4836 2066
rect 4636 1572 4836 1619
rect 4636 1538 4652 1572
rect 4820 1538 4836 1572
rect 4636 1522 4836 1538
<< polycont >>
rect 4552 3186 4720 3220
rect 4552 2658 4720 2692
rect 4652 2066 4820 2100
rect 4652 1538 4820 1572
<< locali >>
rect 4376 3288 4472 3322
rect 4800 3288 4896 3322
rect 4376 3226 4410 3288
rect 4862 3226 4896 3288
rect 4536 3186 4552 3220
rect 4720 3186 4736 3220
rect 4490 3127 4524 3143
rect 4490 2735 4524 2751
rect 4748 3127 4782 3143
rect 4748 2735 4782 2751
rect 4536 2658 4552 2692
rect 4720 2658 4736 2692
rect 4376 2590 4410 2652
rect 4862 2590 4896 2652
rect 4376 2556 4472 2590
rect 4800 2556 4896 2590
rect 4476 2168 4572 2202
rect 4900 2168 4996 2202
rect 4476 2106 4510 2168
rect 4962 2106 4996 2168
rect 4636 2066 4652 2100
rect 4820 2066 4836 2100
rect 4590 2007 4624 2023
rect 4590 1615 4624 1631
rect 4848 2007 4882 2023
rect 4848 1615 4882 1631
rect 4636 1538 4652 1572
rect 4820 1538 4836 1572
rect 4476 1470 4510 1532
rect 4962 1470 4996 1532
rect 4476 1436 4572 1470
rect 4900 1436 4996 1470
<< viali >>
rect 9090 130 9110 210
rect 9110 130 9250 210
rect 9250 130 9270 210
<< metal1 >>
rect 8420 3640 8480 3810
rect 6240 3260 7480 3320
rect 3520 3100 3720 3180
rect 6240 3140 6300 3260
rect 6200 3120 6300 3140
rect 3520 3040 5900 3100
rect 6200 3060 6220 3120
rect 6280 3060 7120 3120
rect 6200 3040 6300 3060
rect 3520 2980 3720 3040
rect 5140 2220 5200 3040
rect 6260 2880 6360 2900
rect 5600 2680 5660 2880
rect 6260 2820 6280 2880
rect 6340 2820 7380 2880
rect 6260 2800 6360 2820
rect 5380 2620 6100 2680
rect 6040 2420 6100 2620
rect 6600 2420 7320 2680
rect 8100 2420 8160 3640
rect 8410 3630 8490 3640
rect 8410 3450 8420 3630
rect 8480 3450 8490 3630
rect 8410 3440 8490 3450
rect 8800 3400 8860 3640
rect 9140 3630 9200 3810
rect 9840 3640 9900 3810
rect 9820 3630 9900 3640
rect 9120 3620 9200 3630
rect 9120 3440 9130 3620
rect 9190 3440 9200 3620
rect 9120 3430 9200 3440
rect 9490 3620 9570 3630
rect 9490 3440 9500 3620
rect 9560 3440 9570 3620
rect 9820 3450 9830 3630
rect 9890 3450 9900 3630
rect 9820 3440 9900 3450
rect 9490 3430 9570 3440
rect 8200 3340 9800 3400
rect 8420 3210 8500 3220
rect 8420 3030 8430 3210
rect 8490 3030 8500 3210
rect 8420 3020 8500 3030
rect 8800 2980 8860 3340
rect 9820 3210 9900 3220
rect 9120 3200 9200 3210
rect 9120 3020 9130 3200
rect 9190 3020 9200 3200
rect 9120 3010 9200 3020
rect 9490 3200 9580 3210
rect 9490 3020 9500 3200
rect 9560 3020 9580 3200
rect 9820 3030 9830 3210
rect 9890 3030 9900 3210
rect 9820 3020 9900 3030
rect 9490 3010 9580 3020
rect 8220 2920 9800 2980
rect 8420 2790 8500 2800
rect 8420 2610 8430 2790
rect 8490 2610 8500 2790
rect 8420 2600 8500 2610
rect 8800 2560 8860 2920
rect 9820 2790 9900 2800
rect 9120 2780 9200 2790
rect 9120 2600 9130 2780
rect 9190 2600 9200 2780
rect 9120 2590 9200 2600
rect 9490 2780 9580 2790
rect 9490 2600 9500 2780
rect 9560 2600 9580 2780
rect 9820 2610 9830 2790
rect 9890 2610 9900 2790
rect 9820 2600 9900 2610
rect 9490 2590 9580 2600
rect 8220 2500 9800 2560
rect 6040 2360 8160 2420
rect 5140 2160 6280 2220
rect 5140 2020 5200 2160
rect 5920 2020 6020 2040
rect 5140 1960 5480 2020
rect 5700 1960 5940 2020
rect 6000 1960 6020 2020
rect 5920 1940 6020 1960
rect 6220 2020 6280 2160
rect 6220 1940 6380 2020
rect 7600 2000 7880 2020
rect 7600 1920 7800 2000
rect 7860 1920 7880 2000
rect 7600 1880 7880 1920
rect 7600 1800 7800 1880
rect 7860 1800 7880 1880
rect 7600 1740 7880 1800
rect 7600 1660 7800 1740
rect 7860 1660 7880 1740
rect 7600 1620 7880 1660
rect 5520 1580 5660 1600
rect 5520 1520 5540 1580
rect 5640 1520 5660 1580
rect 5520 1500 5660 1520
rect 6420 1580 7580 1600
rect 6420 1520 6440 1580
rect 6540 1520 7580 1580
rect 6420 1500 7580 1520
rect 5120 1460 5220 1480
rect 5120 1400 5140 1460
rect 5200 1400 5220 1460
rect 5120 1380 5220 1400
rect 5140 1120 5200 1380
rect 7920 1300 8020 1320
rect 5020 1060 5200 1120
rect 5140 920 5200 1060
rect 3940 860 5200 920
rect 5300 1240 7940 1300
rect 8000 1240 8020 1300
rect 5300 680 5360 1240
rect 7920 1220 8020 1240
rect 7740 1100 7920 1120
rect 7740 1040 7840 1100
rect 7900 1040 7920 1100
rect 7740 1000 7920 1040
rect 7740 940 7840 1000
rect 7900 940 7920 1000
rect 7740 900 7920 940
rect 7740 880 7840 900
rect 5600 840 7840 880
rect 7900 840 7920 900
rect 5600 820 7920 840
rect 4200 620 5360 680
rect 5840 460 7460 680
rect 8100 520 8160 2360
rect 8420 2370 8500 2380
rect 8420 2190 8430 2370
rect 8490 2190 8500 2370
rect 8800 2280 8860 2500
rect 8420 2180 8500 2190
rect 8640 2140 8860 2280
rect 9120 2370 9200 2380
rect 9820 2370 9900 2380
rect 9120 2190 9130 2370
rect 9190 2190 9200 2370
rect 9120 2180 9200 2190
rect 9490 2360 9580 2370
rect 9490 2180 9500 2360
rect 9560 2180 9580 2360
rect 9820 2190 9830 2370
rect 9890 2190 9900 2370
rect 9820 2180 9900 2190
rect 9490 2170 9580 2180
rect 8240 2080 9800 2140
rect 8420 1950 8500 1960
rect 8420 1770 8430 1950
rect 8490 1770 8500 1950
rect 8420 1760 8500 1770
rect 8640 1720 8700 2080
rect 8800 1720 8860 2080
rect 9820 1960 9900 1970
rect 9120 1950 9200 1960
rect 9120 1770 9130 1950
rect 9190 1770 9200 1950
rect 9120 1760 9200 1770
rect 9490 1940 9570 1950
rect 9490 1760 9500 1940
rect 9560 1760 9570 1940
rect 9820 1780 9830 1960
rect 9890 1780 9900 1960
rect 9820 1770 9900 1780
rect 9490 1750 9570 1760
rect 8220 1660 9800 1720
rect 8420 1540 8500 1550
rect 8420 1360 8430 1540
rect 8490 1360 8500 1540
rect 8420 1350 8500 1360
rect 8640 1320 8700 1660
rect 8620 1300 8720 1320
rect 8800 1300 8860 1660
rect 9120 1530 9200 1540
rect 9120 1350 9130 1530
rect 9190 1350 9200 1530
rect 9120 1340 9200 1350
rect 9500 1530 9580 1550
rect 9500 1350 9510 1530
rect 9570 1350 9580 1530
rect 9500 1340 9580 1350
rect 9820 1530 9900 1540
rect 9820 1350 9830 1530
rect 9890 1350 9900 1530
rect 9820 1340 9900 1350
rect 8200 1240 8640 1300
rect 8700 1240 9800 1300
rect 8620 1220 8720 1240
rect 8420 1120 8500 1130
rect 8420 940 8430 1120
rect 8490 940 8500 1120
rect 8420 930 8500 940
rect 8800 900 8860 1240
rect 9120 1120 9200 1130
rect 9120 940 9130 1120
rect 9190 940 9200 1120
rect 9120 920 9200 940
rect 9500 1120 9580 1140
rect 9500 940 9510 1120
rect 9570 940 9580 1120
rect 9500 930 9580 940
rect 9820 1120 9900 1130
rect 9820 940 9830 1120
rect 9890 940 9900 1120
rect 9820 930 9900 940
rect 8200 880 8860 900
rect 8200 840 9800 880
rect 8220 820 9800 840
rect 8420 700 8500 710
rect 8420 520 8430 700
rect 8490 520 8500 700
rect 8420 510 8500 520
rect 8800 480 8860 820
rect 9120 700 9200 710
rect 9120 520 9130 700
rect 9190 520 9200 700
rect 9120 510 9200 520
rect 9500 700 9580 710
rect 9500 520 9510 700
rect 9570 520 9580 700
rect 9500 510 9580 520
rect 9820 700 9900 710
rect 9820 520 9830 700
rect 9890 520 9900 700
rect 9820 510 9900 520
rect 4000 400 7660 460
rect 8180 420 9800 480
rect 5400 380 7660 400
rect 5400 360 9580 380
rect 5400 320 9500 360
rect 5400 240 5600 320
rect 9480 300 9500 320
rect 9560 300 9580 360
rect 9480 280 9580 300
rect 8880 270 9270 280
rect 8880 260 9280 270
rect 5400 160 5420 240
rect 5580 160 5600 240
rect 5400 -60 5600 160
rect 7820 240 7920 260
rect 7820 180 7840 240
rect 7900 180 7920 240
rect 7820 140 7920 180
rect 8880 200 8900 260
rect 9060 210 9280 260
rect 9060 200 9090 210
rect 7760 -60 7960 140
rect 8880 130 9090 200
rect 9270 130 9280 210
rect 8880 110 9280 130
rect 8880 -80 9080 110
<< via1 >>
rect 6220 3060 6280 3120
rect 6280 2820 6340 2880
rect 8420 3450 8480 3630
rect 9130 3440 9190 3620
rect 9500 3440 9560 3620
rect 9830 3450 9890 3630
rect 8430 3030 8490 3210
rect 9130 3020 9190 3200
rect 9500 3020 9560 3200
rect 9830 3030 9890 3210
rect 8430 2610 8490 2790
rect 9130 2600 9190 2780
rect 9500 2600 9560 2780
rect 9830 2610 9890 2790
rect 5940 1960 6000 2020
rect 7800 1920 7860 2000
rect 7800 1800 7860 1880
rect 7800 1660 7860 1740
rect 5540 1520 5640 1580
rect 6440 1520 6540 1580
rect 5140 1400 5200 1460
rect 7940 1240 8000 1300
rect 7840 1040 7900 1100
rect 7840 940 7900 1000
rect 7840 840 7900 900
rect 8430 2190 8490 2370
rect 9130 2190 9190 2370
rect 9500 2180 9560 2360
rect 9830 2190 9890 2370
rect 8430 1770 8490 1950
rect 9130 1770 9190 1950
rect 9500 1760 9560 1940
rect 9830 1780 9890 1960
rect 8430 1360 8490 1540
rect 9130 1350 9190 1530
rect 9510 1350 9570 1530
rect 9830 1350 9890 1530
rect 8640 1240 8700 1300
rect 8430 940 8490 1120
rect 9130 940 9190 1120
rect 9510 940 9570 1120
rect 9830 940 9890 1120
rect 8430 520 8490 700
rect 9130 520 9190 700
rect 9510 520 9570 700
rect 9830 520 9890 700
rect 9500 300 9560 360
rect 5420 160 5580 240
rect 7840 180 7900 240
rect 8900 200 9060 260
<< metal2 >>
rect 8410 3630 8490 3640
rect 9500 3630 9560 3660
rect 9820 3630 9900 3640
rect 8410 3450 8420 3630
rect 8480 3450 8490 3630
rect 8410 3440 8490 3450
rect 9120 3620 9200 3630
rect 9120 3440 9130 3620
rect 9190 3440 9200 3620
rect 9120 3430 9200 3440
rect 9490 3620 9570 3630
rect 9490 3440 9500 3620
rect 9560 3440 9570 3620
rect 9820 3450 9830 3630
rect 9890 3450 9900 3630
rect 9820 3440 9900 3450
rect 9490 3430 9570 3440
rect 8420 3210 8500 3220
rect 9500 3210 9560 3430
rect 9820 3210 9900 3220
rect 6200 3120 6300 3140
rect 5940 3060 6220 3120
rect 6280 3060 6300 3120
rect 5940 2040 6000 3060
rect 6200 3040 6300 3060
rect 8420 3030 8430 3210
rect 8490 3030 8500 3210
rect 8420 3020 8500 3030
rect 9120 3200 9200 3210
rect 9120 3020 9130 3200
rect 9190 3020 9200 3200
rect 9120 3010 9200 3020
rect 9490 3200 9570 3210
rect 9490 3020 9500 3200
rect 9560 3020 9570 3200
rect 9820 3030 9830 3210
rect 9890 3030 9900 3210
rect 9820 3020 9900 3030
rect 9490 3010 9570 3020
rect 6260 2880 6360 2900
rect 6140 2820 6280 2880
rect 6340 2820 6360 2880
rect 5920 2020 6020 2040
rect 5920 1960 5940 2020
rect 6000 1960 6020 2020
rect 5920 1940 6020 1960
rect 5520 1580 5660 1600
rect 5520 1520 5540 1580
rect 5640 1520 5660 1580
rect 5520 1500 5660 1520
rect 5120 1460 5220 1480
rect 6140 1460 6200 2820
rect 6260 2800 6360 2820
rect 8420 2790 8500 2800
rect 9500 2790 9560 3010
rect 9820 2790 9900 2800
rect 8420 2610 8430 2790
rect 8490 2610 8500 2790
rect 8420 2600 8500 2610
rect 9120 2780 9200 2790
rect 9120 2600 9130 2780
rect 9190 2600 9200 2780
rect 9120 2590 9200 2600
rect 9490 2780 9570 2790
rect 9490 2600 9500 2780
rect 9560 2600 9570 2780
rect 9820 2610 9830 2790
rect 9890 2610 9900 2790
rect 9820 2600 9900 2610
rect 9490 2590 9570 2600
rect 8420 2370 8500 2380
rect 8420 2190 8430 2370
rect 8490 2190 8500 2370
rect 8420 2180 8500 2190
rect 9120 2370 9200 2380
rect 9500 2370 9560 2590
rect 9820 2370 9900 2380
rect 9120 2190 9130 2370
rect 9190 2190 9200 2370
rect 9120 2180 9200 2190
rect 9490 2360 9570 2370
rect 9490 2180 9500 2360
rect 9560 2180 9570 2360
rect 9820 2190 9830 2370
rect 9890 2190 9900 2370
rect 9820 2180 9900 2190
rect 9490 2170 9570 2180
rect 7780 2000 7880 2020
rect 7780 1920 7800 2000
rect 7860 1920 7880 2000
rect 7780 1880 7880 1920
rect 7780 1800 7800 1880
rect 7860 1800 7880 1880
rect 7780 1740 7880 1800
rect 8420 1950 8500 1960
rect 8420 1770 8430 1950
rect 8490 1770 8500 1950
rect 8420 1760 8500 1770
rect 9120 1950 9200 1960
rect 9500 1950 9560 2170
rect 9820 1960 9900 1970
rect 9120 1770 9130 1950
rect 9190 1770 9200 1950
rect 9120 1760 9200 1770
rect 9490 1940 9570 1950
rect 9490 1760 9500 1940
rect 9560 1760 9570 1940
rect 9820 1780 9830 1960
rect 9890 1780 9900 1960
rect 9820 1770 9900 1780
rect 9490 1750 9570 1760
rect 7780 1660 7800 1740
rect 7860 1660 7880 1740
rect 7780 1620 7880 1660
rect 6420 1580 6560 1600
rect 6420 1520 6440 1580
rect 6540 1520 6560 1580
rect 6420 1500 6560 1520
rect 5120 1400 5140 1460
rect 5200 1400 6200 1460
rect 5120 1380 5220 1400
rect 7820 1120 7880 1620
rect 8420 1540 8500 1550
rect 9500 1540 9560 1750
rect 8420 1360 8430 1540
rect 8490 1360 8500 1540
rect 8420 1350 8500 1360
rect 9120 1530 9200 1540
rect 9120 1350 9130 1530
rect 9190 1350 9200 1530
rect 9120 1340 9200 1350
rect 9500 1530 9580 1540
rect 9500 1350 9510 1530
rect 9570 1350 9580 1530
rect 9500 1340 9580 1350
rect 9820 1530 9900 1540
rect 9820 1350 9830 1530
rect 9890 1350 9900 1530
rect 9820 1340 9900 1350
rect 7920 1300 8020 1320
rect 8620 1300 8720 1320
rect 7920 1240 7940 1300
rect 8000 1240 8640 1300
rect 8700 1240 8720 1300
rect 7920 1220 8020 1240
rect 8620 1220 8720 1240
rect 9500 1130 9560 1340
rect 8420 1120 8500 1130
rect 7820 1100 7920 1120
rect 7820 1040 7840 1100
rect 7900 1040 7920 1100
rect 7820 1000 7920 1040
rect 7820 940 7840 1000
rect 7900 940 7920 1000
rect 7820 900 7920 940
rect 8420 940 8430 1120
rect 8490 940 8500 1120
rect 8420 930 8500 940
rect 9120 1120 9200 1130
rect 9120 940 9130 1120
rect 9190 940 9200 1120
rect 9120 930 9200 940
rect 9500 1120 9580 1130
rect 9500 940 9510 1120
rect 9570 940 9580 1120
rect 9500 930 9580 940
rect 9820 1120 9900 1130
rect 9820 940 9830 1120
rect 9890 940 9900 1120
rect 9820 930 9900 940
rect 7820 840 7840 900
rect 7900 840 7920 900
rect 7820 820 7920 840
rect 7820 260 7880 820
rect 9500 710 9560 930
rect 8420 700 8500 710
rect 8420 520 8430 700
rect 8490 520 8500 700
rect 8420 510 8500 520
rect 9120 700 9200 710
rect 9120 520 9130 700
rect 9190 520 9200 700
rect 9120 510 9200 520
rect 9500 700 9580 710
rect 9500 520 9510 700
rect 9570 520 9580 700
rect 9500 510 9580 520
rect 9820 700 9900 710
rect 9820 520 9830 700
rect 9890 520 9900 700
rect 9820 510 9900 520
rect 9500 380 9560 510
rect 9480 360 9580 380
rect 9480 300 9500 360
rect 9560 300 9580 360
rect 9480 280 9580 300
rect 8880 260 9080 280
rect 5400 240 5600 260
rect 5400 160 5420 240
rect 5580 160 5600 240
rect 7820 240 7920 260
rect 7820 180 7840 240
rect 7900 180 7920 240
rect 8880 200 8900 260
rect 9060 200 9080 260
rect 8880 180 9080 200
rect 7820 160 7920 180
rect 5400 140 5600 160
<< via2 >>
rect 8420 3450 8480 3630
rect 9130 3440 9190 3620
rect 9830 3450 9890 3630
rect 8430 3030 8490 3210
rect 9130 3020 9190 3200
rect 9830 3030 9890 3210
rect 5540 1520 5640 1580
rect 8430 2610 8490 2790
rect 9130 2600 9190 2780
rect 9830 2610 9890 2790
rect 8430 2190 8490 2370
rect 9130 2190 9190 2370
rect 9830 2190 9890 2370
rect 8430 1770 8490 1950
rect 9130 1770 9190 1950
rect 9830 1780 9890 1960
rect 6440 1520 6540 1580
rect 8430 1360 8490 1540
rect 9130 1350 9190 1530
rect 9830 1350 9890 1530
rect 8430 940 8490 1120
rect 9130 940 9190 1120
rect 9830 940 9890 1120
rect 8430 520 8490 700
rect 9130 520 9190 700
rect 9830 520 9890 700
rect 5420 160 5580 240
rect 8900 200 9060 260
<< metal3 >>
rect 8410 3630 8490 3640
rect 8410 3450 8420 3630
rect 8480 3450 8490 3630
rect 8410 3440 8490 3450
rect 9120 3630 9180 3640
rect 9820 3630 9900 3640
rect 9120 3620 9200 3630
rect 9120 3440 9130 3620
rect 9190 3440 9200 3620
rect 8420 3220 8480 3440
rect 9120 3430 9200 3440
rect 9820 3450 9830 3630
rect 9890 3450 9900 3630
rect 9820 3440 9900 3450
rect 8420 3210 8500 3220
rect 8420 3030 8430 3210
rect 8490 3030 8500 3210
rect 8420 3020 8500 3030
rect 9120 3210 9180 3430
rect 9820 3220 9880 3440
rect 9820 3210 9900 3220
rect 9120 3200 9200 3210
rect 9120 3020 9130 3200
rect 9190 3020 9200 3200
rect 8420 2800 8480 3020
rect 9120 3010 9200 3020
rect 9820 3030 9830 3210
rect 9890 3030 9900 3210
rect 9820 3020 9900 3030
rect 8420 2790 8500 2800
rect 8420 2610 8430 2790
rect 8490 2610 8500 2790
rect 8420 2600 8500 2610
rect 9120 2790 9180 3010
rect 9820 2800 9880 3020
rect 9820 2790 9900 2800
rect 9120 2780 9200 2790
rect 9120 2600 9130 2780
rect 9190 2600 9200 2780
rect 8420 2380 8480 2600
rect 9120 2590 9200 2600
rect 9820 2610 9830 2790
rect 9890 2610 9900 2790
rect 9820 2600 9900 2610
rect 9120 2380 9180 2590
rect 9820 2380 9880 2600
rect 8420 2370 8500 2380
rect 8420 2190 8430 2370
rect 8490 2190 8500 2370
rect 8420 2180 8500 2190
rect 9120 2370 9200 2380
rect 9120 2190 9130 2370
rect 9190 2190 9200 2370
rect 9120 2180 9200 2190
rect 9820 2370 9900 2380
rect 9820 2190 9830 2370
rect 9890 2190 9900 2370
rect 9820 2180 9900 2190
rect 8420 1960 8480 2180
rect 9120 1960 9180 2180
rect 9820 1970 9880 2180
rect 9820 1960 9900 1970
rect 8420 1950 8500 1960
rect 8420 1770 8430 1950
rect 8490 1770 8500 1950
rect 8420 1760 8500 1770
rect 9120 1950 9200 1960
rect 9120 1770 9130 1950
rect 9190 1770 9200 1950
rect 9120 1760 9200 1770
rect 9820 1780 9830 1960
rect 9890 1780 9900 1960
rect 9820 1770 9900 1780
rect 5520 1580 5660 1600
rect 6420 1580 6560 1600
rect 5520 1520 5540 1580
rect 5640 1520 6440 1580
rect 6540 1520 6560 1580
rect 5520 1500 5660 1520
rect 6420 1500 6560 1520
rect 8420 1550 8480 1760
rect 8420 1540 8500 1550
rect 5560 260 5640 1500
rect 5400 240 5640 260
rect 5400 160 5420 240
rect 5580 160 5640 240
rect 8420 1360 8430 1540
rect 8490 1360 8500 1540
rect 8420 1350 8500 1360
rect 9120 1540 9180 1760
rect 9820 1540 9880 1770
rect 9120 1530 9200 1540
rect 9120 1350 9130 1530
rect 9190 1350 9200 1530
rect 8420 1130 8480 1350
rect 9120 1340 9200 1350
rect 9820 1530 9900 1540
rect 9820 1350 9830 1530
rect 9890 1350 9900 1530
rect 9820 1340 9900 1350
rect 9120 1130 9180 1340
rect 9820 1130 9880 1340
rect 8420 1120 8500 1130
rect 8420 940 8430 1120
rect 8490 940 8500 1120
rect 8420 930 8500 940
rect 9120 1120 9200 1130
rect 9120 940 9130 1120
rect 9190 940 9200 1120
rect 8420 710 8480 930
rect 9120 920 9200 940
rect 9820 1120 9900 1130
rect 9820 940 9830 1120
rect 9890 940 9900 1120
rect 9820 930 9900 940
rect 9120 710 9180 920
rect 9820 710 9880 930
rect 8420 700 8500 710
rect 8420 520 8430 700
rect 8490 520 8500 700
rect 8420 510 8500 520
rect 9120 700 9200 710
rect 9120 520 9130 700
rect 9190 520 9200 700
rect 9120 510 9200 520
rect 9820 700 9900 710
rect 9820 520 9830 700
rect 9890 520 9900 700
rect 9820 510 9900 520
rect 8420 280 8480 510
rect 9120 280 9180 510
rect 9820 280 9880 510
rect 8420 260 9880 280
rect 8420 220 8900 260
rect 8880 200 8900 220
rect 9060 220 9880 260
rect 9060 200 9080 220
rect 8880 180 9080 200
rect 5400 140 5640 160
use sky130_fd_pr__nfet_01v8_SXQYJB  XN3
timestamp 1657052488
transform 1 0 9696 0 1 2073
box -296 -1773 296 1773
use sky130_fd_pr__pfet_01v8_8LGM97  XP1
timestamp 1657052488
transform 1 0 5625 0 1 2919
box -425 -419 425 419
use sky130_fd_pr__pfet_01v8_8CLFA7  XP2
timestamp 1657057508
transform 1 0 6954 0 1 2919
box -554 -419 554 419
use sky130_fd_pr__pfet_01v8_G8PMZT  XP3
timestamp 1657052488
transform 1 0 5596 0 1 1819
box -296 -419 296 419
use sky130_fd_pr__pfet_01v8_GA6QLT  XP4
timestamp 1657052488
transform 1 0 6996 0 1 1819
box -796 -419 796 419
use sky130_fd_pr__pfet_01v8_8CL9B7  XP6
timestamp 1657053530
transform 1 0 6647 0 1 701
box -1199 -419 1199 419
use sky130_fd_pr__nfet_01v8_SXQYJB  sky130_fd_pr__nfet_01v8_SXQYJB_0
timestamp 1657052488
transform 1 0 8996 0 1 2073
box -296 -1773 296 1773
use sky130_fd_pr__nfet_01v8_SXQYJB  sky130_fd_pr__nfet_01v8_SXQYJB_1
timestamp 1657052488
transform 1 0 8296 0 1 2073
box -296 -1773 296 1773
use sky130_fd_pr__pfet_01v8_8CLZW6  sky130_fd_pr__pfet_01v8_8CLZW6_0
timestamp 1657052488
transform 1 0 4483 0 1 719
box -683 -419 683 419
<< labels >>
flabel metal1 3520 2980 3720 3180 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 7700 2400 7700 2400 0 FreeSans 800 0 0 0 a
flabel metal2 5960 2360 5960 2360 0 FreeSans 800 0 0 0 d
flabel metal2 6000 1440 6000 1440 0 FreeSans 800 0 0 0 c
flabel metal1 7780 1260 7780 1260 0 FreeSans 800 0 0 0 b
flabel metal1 5400 -60 5600 140 0 FreeSans 1600 0 0 0 vtd
port 2 nsew
flabel metal1 7760 -60 7960 140 0 FreeSans 1600 0 0 0 vts
port 1 nsew
flabel metal1 8880 -80 9080 120 0 FreeSans 1600 0 0 0 gnd
port 3 nsew
<< end >>
