magic
tech sky130A
magscale 1 2
timestamp 1643669011
<< metal1 >>
rect 8800 800 11000 1000
rect 8800 200 9000 800
rect 9600 200 11000 800
rect 8800 0 11000 200
rect 11400 800 13600 1000
rect 11400 200 12800 800
rect 13400 200 13600 800
rect 11400 0 13600 200
rect 4600 -900 5400 -800
rect 4600 -1100 4700 -900
rect 5300 -1100 6700 -900
rect 4600 -1200 5400 -1100
rect 4900 -3400 5100 -1200
rect 10600 -1300 11900 -100
rect 5800 -1500 11900 -1300
rect 5600 -1900 6860 -1780
rect 6100 -3400 6300 -1900
rect 9200 -3400 9400 -1500
rect 13000 -3400 13200 0
<< via1 >>
rect 9000 200 9600 800
rect 12800 200 13400 800
rect 4700 -1100 5300 -900
<< metal2 >>
rect 8800 800 9800 1000
rect 8800 200 9000 800
rect 9600 200 9800 800
rect 8800 0 9800 200
rect 12600 800 13600 1000
rect 12600 200 12800 800
rect 13400 200 13600 800
rect 12600 0 13600 200
rect 4600 -900 5400 -800
rect 4600 -1100 4700 -900
rect 5300 -1100 5400 -900
rect 4600 -1200 5400 -1100
<< via2 >>
rect 9000 200 9600 800
rect 12800 200 13400 800
rect 4700 -1100 5300 -900
<< metal3 >>
rect 13200 6200 14800 6400
rect 13000 2800 14800 6200
rect 13600 1000 14800 2800
rect 8800 800 9800 1000
rect 8800 200 9000 800
rect 9600 200 9800 800
rect 8800 0 9800 200
rect 12600 800 14800 1000
rect 12600 200 12800 800
rect 13400 200 14800 800
rect 12600 0 14800 200
rect 4600 -900 5400 -800
rect 4600 -1100 4700 -900
rect 5300 -1100 5400 -900
rect 4600 -1200 5400 -1100
<< via3 >>
rect 9000 200 9600 800
rect 4700 -1100 5300 -900
<< metal4 >>
rect -2200 33800 25600 34800
rect -2200 6200 -1200 33800
rect -2200 2600 10000 6200
rect -2200 1000 -1200 2600
rect -2200 800 9800 1000
rect -2200 200 9000 800
rect 9600 200 9800 800
rect -2200 0 9800 200
rect 4600 -900 5400 0
rect 4600 -1100 4700 -900
rect 5300 -1100 5400 -900
rect 4600 -1200 5400 -1100
use sky130_fd_pr__nfet_g5v0d10v5_7HVW2G  XM2
timestamp 1643669011
transform 1 0 6245 0 1 -1321
box -844 -678 844 678
use sky130_fd_pr__res_high_po_5p73_2BGFUD  XR0
timestamp 1643669011
transform 0 1 11248 -1 0 539
box -739 -648 739 648
use sky130_fd_pr__cap_mim_m3_1_7KEKME  XC0
timestamp 1643668240
transform 0 1 11275 -1 0 4324
box -2125 -2075 2124 2075
use l0  l0_0
timestamp 1643668240
transform 1 0 -200 0 1 7000
box 0 -1000 27800 27800
<< labels >>
flabel metal1 9200 -3400 9400 -3200 0 FreeSans 256 0 0 0 gnd
port 0 nsew
flabel metal1 6100 -3400 6300 -3200 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 4900 -3400 5100 -3200 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 13000 -3400 13200 -3200 0 FreeSans 256 0 0 0 vd
port 3 nsew
<< end >>
