magic
tech sky130A
magscale 1 2
timestamp 1645729143
<< metal1 >>
rect 8600 -1640 8660 -1620
rect 7700 -1680 9360 -1640
rect 7700 -2760 7720 -1680
rect 8600 -2180 9360 -1680
rect 10360 -1660 11560 -1620
rect 10360 -2100 10960 -1660
rect 11540 -2100 11560 -1660
rect 10360 -2160 11560 -2100
rect 8600 -2760 8680 -2180
rect 8860 -2580 10360 -2240
rect 7700 -2800 8680 -2760
rect 9960 -2800 10360 -2580
rect 6340 -4480 9760 -2800
rect 9880 -3360 10360 -2800
rect 9880 -3740 10660 -3360
rect 9880 -4480 10360 -3740
rect 9718 -4646 9884 -4572
rect 9720 -5160 9880 -4646
rect 6340 -5360 9880 -5160
rect 10480 -5980 10660 -3740
rect 6340 -6180 10660 -5980
rect 10960 -8520 11560 -2160
rect 6340 -9140 11560 -8520
<< via1 >>
rect 7720 -2760 8600 -1680
rect 10960 -2100 11540 -1660
<< metal2 >>
rect 7700 -1680 8660 -1620
rect 7700 -2760 7720 -1680
rect 8600 -2760 8660 -1680
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
rect 7700 -2820 8660 -2760
<< via2 >>
rect 7720 -2760 8600 -1680
rect 10960 -2100 11540 -1660
<< metal3 >>
rect 7700 -1680 8660 -1620
rect 7700 -2760 7720 -1680
rect 8600 -2760 8660 -1680
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
rect 7700 -2820 8660 -2760
<< via3 >>
rect 7720 -2760 8600 -1680
rect 10960 -2100 11540 -1660
<< metal4 >>
rect 7700 -1620 8600 -329
rect 10600 -400 13200 800
rect 12000 -800 13200 -400
rect 7700 -1680 8660 -1620
rect 7700 -2760 7720 -1680
rect 8600 -2760 8660 -1680
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
rect 7700 -2820 8660 -2760
rect 12000 -8800 13200 -1400
<< rmetal4 >>
rect 12000 -1400 13200 -800
<< via4 >>
rect 10960 -2100 11540 -1660
<< metal5 >>
rect 9200 18200 14800 19400
rect 9200 12200 10400 18200
rect 10940 -300 11480 -280
rect 10940 -1600 11580 -300
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
use l0  l0_0
timestamp 1645729143
transform 1 0 -26800 0 1 -50600
box 38800 40000 70000 70000
use sky130_fd_pr__cap_mim_m3_2_QKF9RA  sky130_fd_pr__cap_mim_m3_2_QKF9RA_0
timestamp 1645715600
transform -1 0 9553 0 1 6713
box -2479 -7350 2501 7350
use sky130_fd_pr__nfet_g5v0d10v5_PWYS4E  sky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0
timestamp 1644948032
transform 1 0 9796 0 1 -3646
box -278 -1128 278 1128
use sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN  sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0
timestamp 1644948032
transform 0 1 9872 -1 0 -2093
box -201 -1098 201 1098
<< labels >>
flabel metal1 6340 -3040 6540 -2840 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 6340 -8720 6540 -8520 0 FreeSans 128 0 0 0 vd
port 3 nsew
flabel metal1 6340 -5360 6540 -5160 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 6340 -6180 6540 -5980 0 FreeSans 128 0 0 0 gnd
port 0 nsew
<< end >>
