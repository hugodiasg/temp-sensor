magic
tech sky130A
magscale 1 2
timestamp 1700191285
<< metal1 >>
rect 6000 33780 7320 33820
rect 6000 33500 6940 33780
rect 7260 33500 7320 33780
rect 6000 33480 7320 33500
rect 6040 33140 6240 33480
rect -80 11320 1580 11460
rect 1760 11320 1780 11460
rect -80 11300 1780 11320
rect -320 10720 120 10920
rect 1550 6760 13100 6780
rect 1040 6560 1240 6760
rect 1550 6560 1560 6760
rect 1760 6560 12880 6760
rect 13080 6560 13100 6760
rect 1030 6400 1040 6560
rect 1220 6400 1240 6560
rect 1040 6380 1240 6400
rect 6290 6280 6300 6420
rect 6460 6280 6470 6420
rect 17310 5700 17320 5880
rect 17500 5700 17510 5880
rect 4360 5520 5840 5540
rect 3490 5320 3500 5480
rect 4000 5320 4010 5480
rect 4360 5340 4380 5520
rect 4560 5340 5840 5520
rect 12600 5400 14480 5420
rect 12600 5240 14300 5400
rect 14440 5240 14480 5400
rect 12600 5220 14480 5240
rect 4680 4640 5840 4660
rect 4680 4480 4700 4640
rect 4880 4480 5840 4640
rect 4680 4460 5840 4480
rect 14310 4160 14320 4320
rect 14460 4160 14470 4320
rect 5650 3700 5660 3900
rect 5840 3700 5850 3900
rect 4040 3360 4370 3560
rect 12870 3240 12880 3440
rect 13080 3240 14500 3440
rect 4040 2900 4380 3100
rect 4560 2900 4580 3100
rect 14330 2940 14340 3080
rect 14460 2940 14470 3080
rect 13080 2760 14500 2780
rect 13070 2580 13080 2760
rect 13260 2580 14500 2760
rect 14330 2020 14340 2200
rect 14460 2020 14470 2200
rect 190 40 200 160
rect 480 40 490 160
rect 15830 140 15990 160
rect 14770 0 14930 140
rect 14970 0 15130 140
rect 15230 120 15390 140
rect 15450 120 15610 140
rect 15630 120 15640 140
rect 15190 40 15640 120
rect 15230 0 15390 40
rect 15450 0 15610 40
rect 15630 20 15640 40
rect 15900 120 15990 140
rect 16250 120 16410 140
rect 16450 120 16610 140
rect 15900 40 16610 120
rect 15900 20 15990 40
rect 15650 0 15810 20
rect 16030 -20 16190 40
rect 16250 0 16410 40
rect 16450 0 16610 40
rect 16630 0 16950 140
rect 60 -840 16100 -820
rect 60 -980 200 -840
rect -60 -1140 200 -980
rect 460 -860 16100 -840
rect 460 -880 15680 -860
rect 460 -920 5660 -880
rect 460 -1140 1060 -920
rect -60 -1180 1060 -1140
rect 60 -1200 1060 -1180
rect 1220 -1180 5660 -920
rect 5820 -1100 15680 -880
rect 15880 -1100 16100 -860
rect 5820 -1180 16100 -1100
rect 1220 -1200 16100 -1180
rect 60 -1260 16100 -1200
rect 4680 -1400 4880 -1380
rect 4680 -1500 4700 -1400
rect 4860 -1500 4880 -1400
rect 4680 -1800 4880 -1500
rect 13080 -1400 13280 -1380
rect 13080 -1500 13100 -1400
rect 13260 -1500 13280 -1400
rect 13080 -1800 13280 -1500
rect 14300 -1400 14500 -1380
rect 14300 -1500 14320 -1400
rect 14480 -1500 14500 -1400
rect 14300 -1600 14500 -1500
rect 14280 -1800 14480 -1600
<< via1 >>
rect 6940 33500 7260 33780
rect 1580 11320 1760 11460
rect 1560 6560 1760 6760
rect 12880 6560 13080 6760
rect 1040 6400 1220 6560
rect 6300 6280 6460 6420
rect 17320 5700 17500 5880
rect 3500 5320 4000 5480
rect 4380 5340 4560 5520
rect 14300 5240 14440 5400
rect 4700 4480 4880 4640
rect 14320 4160 14460 4320
rect 5660 3700 5840 3900
rect 12880 3240 13080 3440
rect 4380 2900 4560 3100
rect 14340 2940 14460 3080
rect 13080 2580 13260 2760
rect 14340 2020 14460 2200
rect 200 40 480 160
rect 15640 20 15900 140
rect 200 -1140 460 -840
rect 1060 -1200 1220 -920
rect 5660 -1180 5820 -880
rect 15680 -1100 15880 -860
rect 4700 -1500 4860 -1400
rect 13100 -1500 13260 -1400
rect 14320 -1500 14480 -1400
<< metal2 >>
rect 6940 33780 7260 33790
rect 6940 33490 7260 33500
rect 1560 11460 1780 11500
rect 1560 11320 1580 11460
rect 1760 11320 1780 11460
rect 1560 6760 1780 11320
rect 1040 6560 1220 6570
rect 1760 6560 1780 6760
rect 12880 6760 13100 6780
rect 13080 6560 13100 6760
rect 1560 6550 1760 6560
rect 1040 6390 1220 6400
rect 6300 6420 6460 6430
rect 6300 6270 6460 6280
rect 4360 5520 4560 5540
rect 3500 5480 4000 5490
rect 3500 5310 4000 5320
rect 4360 5340 4380 5520
rect 4360 3100 4560 5340
rect 4360 2900 4380 3100
rect 4380 2890 4560 2900
rect 4660 4640 4880 4680
rect 4660 4480 4700 4640
rect 160 160 500 180
rect 160 40 200 160
rect 480 40 500 160
rect 160 -840 500 40
rect 160 -1140 200 -840
rect 460 -1140 500 -840
rect 160 -1180 500 -1140
rect 1060 -920 1220 -910
rect 1060 -1210 1220 -1200
rect 4660 -1400 4880 4480
rect 5640 3900 5840 3920
rect 5640 3700 5660 3900
rect 5640 -880 5840 3700
rect 12880 3440 13100 6560
rect 17320 5880 17500 5890
rect 17320 5690 17500 5700
rect 14280 5400 14460 5420
rect 14280 5240 14300 5400
rect 14440 5240 14460 5400
rect 14280 4320 14460 5240
rect 14280 4160 14320 4320
rect 14280 4140 14460 4160
rect 13080 3240 13100 3440
rect 12880 3230 13080 3240
rect 14300 3080 14500 3120
rect 14300 2940 14340 3080
rect 14460 2940 14500 3080
rect 5640 -1180 5660 -880
rect 5820 -1180 5840 -880
rect 5640 -1260 5840 -1180
rect 13080 2760 13280 2780
rect 13260 2580 13280 2760
rect 4660 -1500 4700 -1400
rect 4860 -1500 4880 -1400
rect 4660 -1520 4880 -1500
rect 13080 -1400 13280 2580
rect 13080 -1500 13100 -1400
rect 13260 -1500 13280 -1400
rect 13080 -1520 13280 -1500
rect 14300 2200 14500 2940
rect 14300 2020 14340 2200
rect 14460 2020 14500 2200
rect 14300 -1400 14500 2020
rect 15600 140 15940 200
rect 15600 20 15640 140
rect 15900 20 15940 140
rect 15600 -860 15940 20
rect 15600 -1100 15680 -860
rect 15880 -1100 15940 -860
rect 15600 -1180 15940 -1100
rect 14300 -1500 14320 -1400
rect 14480 -1500 14500 -1400
rect 14300 -1520 14500 -1500
<< via2 >>
rect 6940 33500 7260 33780
rect 1040 6400 1220 6560
rect 6300 6280 6460 6420
rect 3500 5320 4000 5480
rect 1060 -1200 1220 -920
rect 17320 5700 17500 5880
<< metal3 >>
rect 6930 33780 7270 33785
rect 6930 33500 6940 33780
rect 7260 33500 7270 33780
rect 6930 33495 7270 33500
rect 1040 6565 1240 6580
rect 1030 6560 1240 6565
rect 1030 6400 1040 6560
rect 1220 6400 1240 6560
rect 6290 6420 6470 6425
rect 1030 6395 1240 6400
rect 1040 -920 1240 6395
rect 6260 6280 6300 6420
rect 6460 6400 7260 6420
rect 6460 6280 6900 6400
rect 7240 6280 7260 6400
rect 6290 6275 6470 6280
rect 6980 5920 17520 5940
rect 6980 5720 7000 5920
rect 7260 5880 17520 5920
rect 7260 5720 17320 5880
rect 6980 5700 17320 5720
rect 17500 5700 17520 5880
rect 17310 5695 17510 5700
rect 3490 5480 4010 5485
rect 3480 5320 3500 5480
rect 4000 5320 6920 5480
rect 3480 5300 6920 5320
rect 7240 5300 7250 5480
rect 3480 5280 7220 5300
rect 1040 -1200 1060 -920
rect 1220 -1200 1240 -920
rect 1040 -1260 1240 -1200
<< via3 >>
rect 6940 33500 7260 33780
rect 6900 6280 7240 6400
rect 7000 5720 7260 5920
rect 6920 5300 7240 5480
<< metal4 >>
rect 6900 33780 7280 33860
rect 6900 33500 6940 33780
rect 7260 33500 7280 33780
rect 6900 6401 7280 33500
rect 6899 6400 7280 6401
rect 6899 6280 6900 6400
rect 7240 6280 7280 6400
rect 6899 6279 7280 6280
rect 6900 5920 7280 6279
rect 6900 5720 7000 5920
rect 7260 5720 7280 5920
rect 6900 5480 7280 5720
rect 6900 5300 6920 5480
rect 7240 5300 7280 5480
rect 6900 5150 7280 5300
use ask-modulator  ask-modulator_0 /foss/designs/temp-sensor/ask_modulator/mag
timestamp 1700191285
transform 1 0 -740 0 1 16920
box 660 -10360 23078 16420
use buffer  buffer_0 /foss/designs/temp-sensor/buffer/mag
timestamp 1700177945
transform 1 0 -4120 0 1 2820
box 9760 -2860 16933 3620
use sensor  sensor_0 /foss/designs/temp-sensor/sensor/mag
timestamp 1699935153
transform 1 0 660 0 1 2500
box -660 -2500 3580 3000
use sigma-delta  sigma-delta_0 /foss/designs/temp-sensor/sigma-delta_modulator/mag
timestamp 1700102200
transform 1 0 17480 0 1 520
box -3180 -520 5760 5360
<< labels >>
flabel metal1 6040 33620 6240 33820 0 FreeSans 6400 0 0 0 vd
port 0 nsew
flabel metal1 -60 -1180 140 -980 0 FreeSans 6400 0 0 0 gnd
port 1 nsew
flabel metal1 -320 10720 -120 10920 0 FreeSans 6400 0 0 0 out
port 3 nsew
flabel metal1 4680 -1800 4880 -1600 0 FreeSans 6400 0 0 0 ib
port 5 nsew
flabel metal1 14280 -1800 14480 -1600 0 FreeSans 6400 0 0 0 vpwr
port 4 nsew
flabel metal1 13080 -1800 13280 -1600 0 FreeSans 6400 0 0 0 clk
port 2 nsew
flabel metal1 5262 5516 5292 5520 0 FreeSans 1600 0 0 0 vts
flabel metal1 4306 3508 4334 3538 0 FreeSans 1600 0 0 0 vtd
flabel metal1 13376 5282 13494 5370 0 FreeSans 1600 0 0 0 out_buff
flabel metal1 11842 6654 11886 6698 0 FreeSans 800 0 0 0 out_sigma
<< end >>
