magic
tech sky130A
magscale 1 2
timestamp 1645644904
<< metal4 >>
rect -2679 7859 2679 7900
rect -2679 2741 2423 7859
rect 2659 2741 2679 7859
rect -2679 2700 2679 2741
rect -2679 2559 2679 2600
rect -2679 -2559 2423 2559
rect 2659 -2559 2679 2559
rect -2679 -2600 2679 -2559
rect -2679 -2741 2679 -2700
rect -2679 -7859 2423 -2741
rect 2659 -7859 2679 -2741
rect -2679 -7900 2679 -7859
<< via4 >>
rect 2423 2741 2659 7859
rect 2423 -2559 2659 2559
rect 2423 -7859 2659 -2741
<< mimcap2 >>
rect -2579 7760 2421 7800
rect -2579 2840 -2047 7760
rect 1889 2840 2421 7760
rect -2579 2800 2421 2840
rect -2579 2460 2421 2500
rect -2579 -2460 -2047 2460
rect 1889 -2460 2421 2460
rect -2579 -2500 2421 -2460
rect -2579 -2840 2421 -2800
rect -2579 -7760 -2047 -2840
rect 1889 -7760 2421 -2840
rect -2579 -7800 2421 -7760
<< mimcap2contact >>
rect -2047 2840 1889 7760
rect -2047 -2460 1889 2460
rect -2047 -7760 1889 -2840
<< metal5 >>
rect -239 7784 81 7950
rect 2381 7859 2701 7950
rect -2071 7760 1913 7784
rect -2071 2840 -2047 7760
rect 1889 2840 1913 7760
rect -2071 2816 1913 2840
rect -239 2484 81 2816
rect 2381 2741 2423 7859
rect 2659 2741 2701 7859
rect 2381 2559 2701 2741
rect -2071 2460 1913 2484
rect -2071 -2460 -2047 2460
rect 1889 -2460 1913 2460
rect -2071 -2484 1913 -2460
rect -239 -2816 81 -2484
rect 2381 -2559 2423 2559
rect 2659 -2559 2701 2559
rect 2381 -2741 2701 -2559
rect -2071 -2840 1913 -2816
rect -2071 -7760 -2047 -2840
rect 1889 -7760 1913 -2840
rect -2071 -7784 1913 -7760
rect -239 -7950 81 -7784
rect 2381 -7859 2423 -2741
rect 2659 -7859 2701 -2741
rect 2381 -7950 2701 -7859
<< properties >>
string FIXED_BBOX -2679 2700 2521 7900
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25 l 25 val 1.269k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
