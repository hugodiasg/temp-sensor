magic
tech sky130A
magscale 1 2
timestamp 1644768117
<< metal4 >>
rect -2529 7409 2529 7450
rect -2529 2591 2273 7409
rect 2509 2591 2529 7409
rect -2529 2550 2529 2591
rect -2529 2409 2529 2450
rect -2529 -2409 2273 2409
rect 2509 -2409 2529 2409
rect -2529 -2450 2529 -2409
rect -2529 -2591 2529 -2550
rect -2529 -7409 2273 -2591
rect 2509 -7409 2529 -2591
rect -2529 -7450 2529 -7409
<< via4 >>
rect 2273 2591 2509 7409
rect 2273 -2409 2509 2409
rect 2273 -7409 2509 -2591
<< mimcap2 >>
rect -2429 7310 2271 7350
rect -2429 2690 -1927 7310
rect 1769 2690 2271 7310
rect -2429 2650 2271 2690
rect -2429 2310 2271 2350
rect -2429 -2310 -1927 2310
rect 1769 -2310 2271 2310
rect -2429 -2350 2271 -2310
rect -2429 -2690 2271 -2650
rect -2429 -7310 -1927 -2690
rect 1769 -7310 2271 -2690
rect -2429 -7350 2271 -7310
<< mimcap2contact >>
rect -1927 2690 1769 7310
rect -1927 -2310 1769 2310
rect -1927 -7310 1769 -2690
<< metal5 >>
rect -239 7334 81 7500
rect 2231 7409 2551 7500
rect -1951 7310 1793 7334
rect -1951 2690 -1927 7310
rect 1769 2690 1793 7310
rect -1951 2666 1793 2690
rect -239 2334 81 2666
rect 2231 2591 2273 7409
rect 2509 2591 2551 7409
rect 2231 2409 2551 2591
rect -1951 2310 1793 2334
rect -1951 -2310 -1927 2310
rect 1769 -2310 1793 2310
rect -1951 -2334 1793 -2310
rect -239 -2666 81 -2334
rect 2231 -2409 2273 2409
rect 2509 -2409 2551 2409
rect 2231 -2591 2551 -2409
rect -1951 -2690 1793 -2666
rect -1951 -7310 -1927 -2690
rect 1769 -7310 1793 -2690
rect -1951 -7334 1793 -7310
rect -239 -7500 81 -7334
rect 2231 -7409 2273 -2591
rect 2509 -7409 2551 -2591
rect 2231 -7500 2551 -7409
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2529 2550 2371 7450
string parameters w 23.5 l 23.5 val 1.122k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
