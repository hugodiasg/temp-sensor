magic
tech sky130A
magscale 1 2
timestamp 1646100680
<< metal4 >>
rect -2619 10269 2619 10310
rect -2619 5271 2363 10269
rect 2599 5271 2619 10269
rect -2619 5230 2619 5271
rect -2619 5089 2619 5130
rect -2619 91 2363 5089
rect 2599 91 2619 5089
rect -2619 50 2619 91
rect -2619 -91 2619 -50
rect -2619 -5089 2363 -91
rect 2599 -5089 2619 -91
rect -2619 -5130 2619 -5089
rect -2619 -5271 2619 -5230
rect -2619 -10269 2363 -5271
rect 2599 -10269 2619 -5271
rect -2619 -10310 2619 -10269
<< via4 >>
rect 2363 5271 2599 10269
rect 2363 91 2599 5089
rect 2363 -5089 2599 -91
rect 2363 -10269 2599 -5271
<< mimcap2 >>
rect -2519 10170 2361 10210
rect -2519 5370 -1999 10170
rect 1841 5370 2361 10170
rect -2519 5330 2361 5370
rect -2519 4990 2361 5030
rect -2519 190 -1999 4990
rect 1841 190 2361 4990
rect -2519 150 2361 190
rect -2519 -190 2361 -150
rect -2519 -4990 -1999 -190
rect 1841 -4990 2361 -190
rect -2519 -5030 2361 -4990
rect -2519 -5370 2361 -5330
rect -2519 -10170 -1999 -5370
rect 1841 -10170 2361 -5370
rect -2519 -10210 2361 -10170
<< mimcap2contact >>
rect -1999 5370 1841 10170
rect -1999 190 1841 4990
rect -1999 -4990 1841 -190
rect -1999 -10170 1841 -5370
<< metal5 >>
rect -239 10194 81 10360
rect 2321 10269 2641 10360
rect -2023 10170 1865 10194
rect -2023 5370 -1999 10170
rect 1841 5370 1865 10170
rect -2023 5346 1865 5370
rect -239 5014 81 5346
rect 2321 5271 2363 10269
rect 2599 5271 2641 10269
rect 2321 5089 2641 5271
rect -2023 4990 1865 5014
rect -2023 190 -1999 4990
rect 1841 190 1865 4990
rect -2023 166 1865 190
rect -239 -166 81 166
rect 2321 91 2363 5089
rect 2599 91 2641 5089
rect 2321 -91 2641 91
rect -2023 -190 1865 -166
rect -2023 -4990 -1999 -190
rect 1841 -4990 1865 -190
rect -2023 -5014 1865 -4990
rect -239 -5346 81 -5014
rect 2321 -5089 2363 -91
rect 2599 -5089 2641 -91
rect 2321 -5271 2641 -5089
rect -2023 -5370 1865 -5346
rect -2023 -10170 -1999 -5370
rect 1841 -10170 1865 -5370
rect -2023 -10194 1865 -10170
rect -239 -10360 81 -10194
rect 2321 -10269 2363 -5271
rect 2599 -10269 2641 -5271
rect 2321 -10360 2641 -10269
<< properties >>
string FIXED_BBOX -2619 5230 2461 10310
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.399 l 24.399 val 1.209k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
