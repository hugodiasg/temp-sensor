magic
tech sky130A
magscale 1 2
timestamp 1644359060
<< metal1 >>
rect 15736 8200 16200 8858
rect 15700 7300 16200 8200
rect 11800 7200 16200 7300
rect 11800 6400 11900 7200
rect 12700 6400 16200 7200
rect 11800 6200 16200 6400
rect 14980 2760 15380 6200
rect 15675 5200 16200 6200
rect 16500 7300 17200 8900
rect 16500 7200 20700 7300
rect 16500 6400 19800 7200
rect 20600 6400 20700 7200
rect 16500 6200 20700 6400
rect 15675 4994 16043 5200
rect 16500 5000 17200 6200
rect 15675 4732 17186 4843
rect 15675 4676 17180 4732
rect 15669 4525 17180 4676
rect 15669 4096 17164 4525
rect 17337 4096 17480 4100
rect 15669 3505 17480 4096
rect 15700 3500 17480 3505
rect 16700 3200 17480 3500
rect 14980 1980 16320 2760
rect 16440 2600 17480 3200
rect 14980 -320 15380 1980
rect 16200 -320 16600 1620
rect 17080 1163 17480 2600
rect 17080 867 17477 1163
rect 17080 -311 17486 867
rect 17080 -320 17480 -311
rect 18700 -320 19100 6200
rect 15080 -520 15280 -320
rect 16300 -520 16500 -320
rect 17160 -520 17360 -320
rect 18800 -520 19000 -320
<< via1 >>
rect 11900 6400 12700 7200
rect 19800 6400 20600 7200
<< metal2 >>
rect 11800 7200 12800 7300
rect 11800 6400 11900 7200
rect 12700 6400 12800 7200
rect 11800 6200 12800 6400
rect 19700 7200 20700 7300
rect 19700 6400 19800 7200
rect 20600 6400 20700 7200
rect 19700 6200 20700 6400
<< via2 >>
rect 11900 6400 12700 7200
rect 19800 6400 20600 7200
<< metal3 >>
rect 11800 7200 12800 7300
rect 11800 6400 11900 7200
rect 12700 6400 12800 7200
rect 11800 6200 12800 6400
rect 19700 7200 20700 7300
rect 19700 6400 19800 7200
rect 20600 6400 20700 7200
rect 19700 6200 20700 6400
<< via3 >>
rect 11900 6400 12700 7200
rect 19800 6400 20600 7200
<< metal4 >>
rect 11800 27100 39100 28100
rect 11800 7200 12800 27100
rect 16200 24100 17100 27100
rect 38100 19100 39100 27100
rect 11800 6400 11900 7200
rect 12700 6400 12800 7200
rect 11800 6200 12800 6400
rect 19700 7200 20700 7300
rect 19700 6400 19800 7200
rect 20600 6400 20700 7200
rect 19700 6200 20700 6400
<< via4 >>
rect 30100 19200 30900 20000
rect 19800 6400 20600 7200
<< metal5 >>
rect 16200 25500 34900 26500
rect 16200 24100 17100 25500
rect 19700 7200 20700 25500
rect 30076 20000 30924 20024
rect 30076 19200 30100 20000
rect 30900 19200 30924 20000
rect 30076 19176 30924 19200
rect 19700 6400 19800 7200
rect 20600 6400 20700 7200
rect 19700 6200 20700 6400
use l0  l0_0
timestamp 1644072167
transform 1 0 21200 0 1 10300
box 0 0 17200 16200
use sky130_fd_pr__cap_mim_m3_2_QKF9RA  sky130_fd_pr__cap_mim_m3_2_QKF9RA_0
timestamp 1644357294
transform 1 0 16479 0 1 17030
box -2479 -7350 2501 7350
use sky130_fd_pr__res_high_po_5p73_K9JT5B  XR0
timestamp 1644357294
transform 0 1 16446 -1 0 6898
box -2133 -654 2133 654
use sky130_fd_pr__nfet_g5v0d10v5_FLFTBY  XM2
timestamp 1644164861
transform -1 0 16398 0 1 2488
box -278 -1128 278 1128
<< labels >>
flabel metal1 17160 -520 17360 -320 0 FreeSans 128 0 0 0 gnd
port 0 nsew
flabel metal1 18800 -520 19000 -320 0 FreeSans 128 0 0 0 vd
port 3 nsew
flabel metal1 15080 -520 15280 -320 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 16300 -520 16500 -320 0 FreeSans 128 0 0 0 in
port 1 nsew
<< end >>
