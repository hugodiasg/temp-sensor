** sch_path: /home/hugodg/projects-sky130/temp-sensor/sensor/xschem/sensor.sch
.subckt sensor vd vts vtd gnd
*.PININFO vd:B vts:O vtd:O gnd:B
XP1 a a vd vd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=2 m=1
XP2 c a d d sky130_fd_pr__pfet_01v8 L=1 W=8 nf=4 m=1
XP3 d vtd vd vd sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XP4 vts vtd vd vd sky130_fd_pr__pfet_01v8 L=5 W=2 nf=1 m=1
XP5 b vtd c c sky130_fd_pr__pfet_01v8 L=1 W=8 nf=4 m=1
XP6 vtd vtd vts vts sky130_fd_pr__pfet_01v8 L=1 W=16 nf=8 m=1
XN1 a b gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=8
XN2 b b gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=8
XN3 vtd b gnd gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=8
XPD1 net4 net1 net3 net2 sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XPD2 net8 net5 net7 net6 sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XPD3 net12 net9 net11 net10 sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XPD4 net16 net13 net15 net14 sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XPD5 net20 net17 net19 net18 sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XND1 net22 net21 net23 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND2 net25 net24 net26 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND3 net28 net27 net29 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND4 net31 net30 net32 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND5 net34 net33 net35 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND6 net37 net36 net38 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND7 net40 net39 net41 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XND8 net43 net42 net44 gnd sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
.ends
.end
