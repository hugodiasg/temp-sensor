magic
tech sky130A
magscale 1 2
timestamp 1675569099
<< metal4 >>
rect -2669 22519 2669 22560
rect -2669 17801 2413 22519
rect 2649 17801 2669 22519
rect -2669 17760 2669 17801
rect -2669 17479 2669 17520
rect -2669 12761 2413 17479
rect 2649 12761 2669 17479
rect -2669 12720 2669 12761
rect -2669 12439 2669 12480
rect -2669 7721 2413 12439
rect 2649 7721 2669 12439
rect -2669 7680 2669 7721
rect -2669 7399 2669 7440
rect -2669 2681 2413 7399
rect 2649 2681 2669 7399
rect -2669 2640 2669 2681
rect -2669 2359 2669 2400
rect -2669 -2359 2413 2359
rect 2649 -2359 2669 2359
rect -2669 -2400 2669 -2359
rect -2669 -2681 2669 -2640
rect -2669 -7399 2413 -2681
rect 2649 -7399 2669 -2681
rect -2669 -7440 2669 -7399
rect -2669 -7721 2669 -7680
rect -2669 -12439 2413 -7721
rect 2649 -12439 2669 -7721
rect -2669 -12480 2669 -12439
rect -2669 -12761 2669 -12720
rect -2669 -17479 2413 -12761
rect 2649 -17479 2669 -12761
rect -2669 -17520 2669 -17479
rect -2669 -17801 2669 -17760
rect -2669 -22519 2413 -17801
rect 2649 -22519 2669 -17801
rect -2669 -22560 2669 -22519
<< via4 >>
rect 2413 17801 2649 22519
rect 2413 12761 2649 17479
rect 2413 7721 2649 12439
rect 2413 2681 2649 7399
rect 2413 -2359 2649 2359
rect 2413 -7399 2649 -2681
rect 2413 -12439 2649 -7721
rect 2413 -17479 2649 -12761
rect 2413 -22519 2649 -17801
<< mimcap2 >>
rect -2589 22440 2051 22480
rect -2589 17880 -2549 22440
rect 2011 17880 2051 22440
rect -2589 17840 2051 17880
rect -2589 17400 2051 17440
rect -2589 12840 -2549 17400
rect 2011 12840 2051 17400
rect -2589 12800 2051 12840
rect -2589 12360 2051 12400
rect -2589 7800 -2549 12360
rect 2011 7800 2051 12360
rect -2589 7760 2051 7800
rect -2589 7320 2051 7360
rect -2589 2760 -2549 7320
rect 2011 2760 2051 7320
rect -2589 2720 2051 2760
rect -2589 2280 2051 2320
rect -2589 -2280 -2549 2280
rect 2011 -2280 2051 2280
rect -2589 -2320 2051 -2280
rect -2589 -2760 2051 -2720
rect -2589 -7320 -2549 -2760
rect 2011 -7320 2051 -2760
rect -2589 -7360 2051 -7320
rect -2589 -7800 2051 -7760
rect -2589 -12360 -2549 -7800
rect 2011 -12360 2051 -7800
rect -2589 -12400 2051 -12360
rect -2589 -12840 2051 -12800
rect -2589 -17400 -2549 -12840
rect 2011 -17400 2051 -12840
rect -2589 -17440 2051 -17400
rect -2589 -17880 2051 -17840
rect -2589 -22440 -2549 -17880
rect 2011 -22440 2051 -17880
rect -2589 -22480 2051 -22440
<< mimcap2contact >>
rect -2549 17880 2011 22440
rect -2549 12840 2011 17400
rect -2549 7800 2011 12360
rect -2549 2760 2011 7320
rect -2549 -2280 2011 2280
rect -2549 -7320 2011 -2760
rect -2549 -12360 2011 -7800
rect -2549 -17400 2011 -12840
rect -2549 -22440 2011 -17880
<< metal5 >>
rect -429 22464 -109 22680
rect 2371 22519 2691 22680
rect -2573 22440 2035 22464
rect -2573 17880 -2549 22440
rect 2011 17880 2035 22440
rect -2573 17856 2035 17880
rect -429 17424 -109 17856
rect 2371 17801 2413 22519
rect 2649 17801 2691 22519
rect 2371 17479 2691 17801
rect -2573 17400 2035 17424
rect -2573 12840 -2549 17400
rect 2011 12840 2035 17400
rect -2573 12816 2035 12840
rect -429 12384 -109 12816
rect 2371 12761 2413 17479
rect 2649 12761 2691 17479
rect 2371 12439 2691 12761
rect -2573 12360 2035 12384
rect -2573 7800 -2549 12360
rect 2011 7800 2035 12360
rect -2573 7776 2035 7800
rect -429 7344 -109 7776
rect 2371 7721 2413 12439
rect 2649 7721 2691 12439
rect 2371 7399 2691 7721
rect -2573 7320 2035 7344
rect -2573 2760 -2549 7320
rect 2011 2760 2035 7320
rect -2573 2736 2035 2760
rect -429 2304 -109 2736
rect 2371 2681 2413 7399
rect 2649 2681 2691 7399
rect 2371 2359 2691 2681
rect -2573 2280 2035 2304
rect -2573 -2280 -2549 2280
rect 2011 -2280 2035 2280
rect -2573 -2304 2035 -2280
rect -429 -2736 -109 -2304
rect 2371 -2359 2413 2359
rect 2649 -2359 2691 2359
rect 2371 -2681 2691 -2359
rect -2573 -2760 2035 -2736
rect -2573 -7320 -2549 -2760
rect 2011 -7320 2035 -2760
rect -2573 -7344 2035 -7320
rect -429 -7776 -109 -7344
rect 2371 -7399 2413 -2681
rect 2649 -7399 2691 -2681
rect 2371 -7721 2691 -7399
rect -2573 -7800 2035 -7776
rect -2573 -12360 -2549 -7800
rect 2011 -12360 2035 -7800
rect -2573 -12384 2035 -12360
rect -429 -12816 -109 -12384
rect 2371 -12439 2413 -7721
rect 2649 -12439 2691 -7721
rect 2371 -12761 2691 -12439
rect -2573 -12840 2035 -12816
rect -2573 -17400 -2549 -12840
rect 2011 -17400 2035 -12840
rect -2573 -17424 2035 -17400
rect -429 -17856 -109 -17424
rect 2371 -17479 2413 -12761
rect 2649 -17479 2691 -12761
rect 2371 -17801 2691 -17479
rect -2573 -17880 2035 -17856
rect -2573 -22440 -2549 -17880
rect 2011 -22440 2035 -17880
rect -2573 -22464 2035 -22440
rect -429 -22680 -109 -22464
rect 2371 -22519 2413 -17801
rect 2649 -22519 2691 -17801
rect 2371 -22680 2691 -22519
<< properties >>
string FIXED_BBOX -2669 17760 2131 22560
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.2 l 23.2 val 1.094k carea 2.00 cperi 0.19 nx 1 ny 9 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
