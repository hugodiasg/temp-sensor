* NGSPICE file created from device-complete.ext - technology: sky130A

.subckt sensor vd vts vtd gnd
X0 b vtd c vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X1 gnd b b gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 vtd b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 vtd b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=11.6 ps=103 w=1 l=1
X5 vts vtd vtd vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 gnd b vtd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X7 gnd b vtd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X8 vts vtd vtd vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X9 gnd b b gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X10 gnd b b gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 c vtd b vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X12 vtd vtd vts vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 gnd b a gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X14 d vtd vd vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X15 c vtd b vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 b b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X17 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X18 b b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X19 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X20 a a vd vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X21 a b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X22 a b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X23 vd a a vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X24 vtd b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X25 vts vtd vtd vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X27 vd vd vd vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=5.22 ps=41.2 w=2 l=1
X28 b vtd c vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 vtd b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X30 gnd b vtd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X31 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X32 c a d vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X33 vtd vtd vts vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X35 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X36 vd vd vd vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X37 d a c vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X38 b b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X39 gnd b b gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X40 vd vd vd vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X41 c a d vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X42 vtd vtd vts vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X43 gnd b a gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X44 d a c vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X45 gnd b a gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X46 gnd b a gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X47 b b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X48 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X49 gnd b vtd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X50 a b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X51 vts vts vts vts sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=5.22 ps=41.2 w=2 l=1
X52 vts vtd vtd vts sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X53 vd vtd vts vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X54 vtd vtd vts vts sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X55 c c c vd sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=1
X56 vts vts vts vts sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X57 a b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt buffer vd ib out in gnd
X0 b b vd vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 vd vd vd vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=11 ps=81.8 w=1 l=1
X2 c out a gnd sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X3 out d gnd gnd sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a a a vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=1.16 ps=10.3 w=1 l=1
X5 d a vd vd sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X6 d d d vd sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=17.4 ps=122 w=15 l=1
X7 vd vd vd vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X8 a a vd vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X9 gnd d out gnd sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 vd b out vd sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X11 out out out vd sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=17.4 ps=122 w=15 l=1
X12 d d gnd gnd sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a a vd vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 b b b vd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=1.16 ps=10.3 w=1 l=1
X15 a a a gnd sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0.96 ps=7.28 w=1.5 l=0.15
X16 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=7.54 ps=55.5 w=5 l=1
X17 vd a a vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X18 vd a a vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X19 a a vd vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 b b b gnd sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.96 ps=7.28 w=1.5 l=0.15
X21 gnd ib ib gnd sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 c ib gnd gnd sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 ib ib ib gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.58 ps=5.16 w=1 l=1
X24 out b vd vd sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X25 b b vd vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 vd b b vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 gnd d d gnd sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 out out out vd sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0 w=15 l=1
X29 vd b b vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X30 b in c gnd sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X31 c c c gnd sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=1.08 ps=8.82 w=1 l=1
X32 vd a d vd sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X33 d d d vd sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0 w=15 l=1
X34 out d sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X35 vd b b vd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=1
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_7RFGLT a_n165_n1062# a_n35_500# a_n35_n932#
X0 a_n35_500# a_n35_n932# a_n165_n1062# sky130_fd_pr__res_xhigh_po_0p35 l=5
.ends

.subckt sky130_fd_pr__nfet_01v8_LPSAWK a_15_n200# a_n175_n374# a_n73_n200# a_n33_n288#
X0 a_15_n200# a_n33_n288# a_n73_n200# a_n175_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_5FNSJ7 m4_n2789_n7800# c2_n2709_n7720#
X0 c2_n2709_n7720# m4_n2789_n7800# sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X1 c2_n2709_n7720# m4_n2789_n7800# sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X2 c2_n2709_n7720# m4_n2789_n7800# sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
.ends

.subckt ask-modulator in out vd gnd
XXR1 gnd vd out sky130_fd_pr__res_xhigh_po_0p35_7RFGLT
XXM1 gnd gnd out in sky130_fd_pr__nfet_01v8_LPSAWK
XXC0 out vd sky130_fd_pr__cap_mim_m3_2_5FNSJ7
.ends

.subckt sigma-delta gnd vd in a_n3084_1636# x1/VGND clk out reset_b_dff vpwr
X0 a_n1599_309# a_n1774_335# a_n1420_335# gnd sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1 a_n2266_4800# a_n2100_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X2 a_n1124_4800# a_n958_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X3 x1.Q a_n1599_309# vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.213 ps=1.67 w=1 l=0.15
X4 a_n2339_335# a_n2689_335# a_n2434_335# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5 a_n2121_577# a_n2339_335# vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X6 a_n1420_335# reset_b_dff gnd gnd sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X7 a_n792_4800# a_n626_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X8 in_int gnd sky130_fd_pr__cap_mim_m3_2 l=27.2 w=27.2
X9 a_n2714_2632# a_n2880_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X10 out a_n1035_335# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X11 a_n1934_4800# a_n2100_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X12 in_comp a_n1884_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X13 a_n1612_701# a_n2689_335# a_n1774_335# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 a_n2077_335# a_n2121_577# a_n2243_335# gnd sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X15 a_n2434_335# x1.D gnd gnd sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 a_n1599_309# reset_b_dff vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X17 a_n2598_4800# a_n2764_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X18 a_n1665_335# a_n2855_335# a_n1774_335# gnd sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X19 a_n1456_4800# in_int gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X20 gnd a_n1599_309# a_n1665_335# gnd sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X21 a_n2434_335# x1.D vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X22 vpwr a_n1599_309# a_n1612_701# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 vpwr a_n1774_335# a_n1599_309# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 a_n2121_577# a_n2339_335# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X25 vpwr clk a_n2855_335# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X26 gnd reset_b_dff a_n2077_335# gnd sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X27 vpwr a_n1599_309# a_n1035_335# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X28 gnd a_n1599_309# a_n1035_335# gnd sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_n2266_4800# a_n2432_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X30 a_n2050_2632# a_n2216_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X31 gnd clk a_n2855_335# gnd sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_n2243_335# a_n2689_335# a_n2339_335# gnd sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X33 vd in_comp x1.D vd sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X34 a_n1124_4800# a_n1290_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X35 a_n2339_335# a_n2855_335# a_n2434_335# gnd sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X36 a_n460_4800# x1.Q gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X37 a_n2689_335# a_n2855_335# vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X38 a_n2231_701# a_n2855_335# a_n2339_335# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X39 a_n2689_335# a_n2855_335# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X40 a_n1774_335# a_n2855_335# a_n2121_577# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X41 a_n2382_2632# a_n2548_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X42 in_int a_n2880_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X43 x1.Q a_n1599_309# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X44 a_n460_4800# a_n626_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X45 a_n2231_701# reset_b_dff vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X46 a_n2930_4800# a_n2764_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X47 a_n2714_2632# a_n2548_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X48 gnd in_comp x1.D gnd sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X49 a_n1934_4800# in_int gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X50 a_n792_4800# a_n958_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X51 vpwr a_n2121_577# a_n2231_701# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X52 a_n1774_335# a_n2689_335# a_n2121_577# gnd sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X53 a_n2598_4800# a_n2432_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X54 a_n2382_2632# a_n2216_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X55 in_comp gnd sky130_fd_pr__cap_mim_m3_2 l=27.2 w=27.2
X56 a_n2930_4800# in gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X57 a_n1456_4800# a_n1290_3468# gnd sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X58 a_n2050_2632# a_n1884_1800# gnd sky130_fd_pr__res_xhigh_po_0p35 l=2
X59 out a_n1035_335# vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
.ends

.subckt device-complete vd gnd clk out vpwr ib out_buff vts out_sigma
Xsensor_0 vd vts vtd gnd sensor
Xbuffer_0 vd ib out_buff vts gnd buffer
Xask-modulator_0 out_sigma out vd gnd ask-modulator
Xsigma-delta_0 gnd vd out_buff gnd gnd clk out_sigma vpwr vpwr sigma-delta
.ends

