magic
tech sky130A
magscale 1 2
timestamp 1645800166
<< metal4 >>
rect -2675 10493 2675 10534
rect -2675 5383 2419 10493
rect 2655 5383 2675 10493
rect -2675 5342 2675 5383
rect -2675 5201 2675 5242
rect -2675 91 2419 5201
rect 2655 91 2675 5201
rect -2675 50 2675 91
rect -2675 -91 2675 -50
rect -2675 -5201 2419 -91
rect 2655 -5201 2675 -91
rect -2675 -5242 2675 -5201
rect -2675 -5383 2675 -5342
rect -2675 -10493 2419 -5383
rect 2655 -10493 2675 -5383
rect -2675 -10534 2675 -10493
<< via4 >>
rect 2419 5383 2655 10493
rect 2419 91 2655 5201
rect 2419 -5201 2655 -91
rect 2419 -10493 2655 -5383
<< mimcap2 >>
rect -2575 10394 2417 10434
rect -2575 5482 -2044 10394
rect 1886 5482 2417 10394
rect -2575 5442 2417 5482
rect -2575 5102 2417 5142
rect -2575 190 -2044 5102
rect 1886 190 2417 5102
rect -2575 150 2417 190
rect -2575 -190 2417 -150
rect -2575 -5102 -2044 -190
rect 1886 -5102 2417 -190
rect -2575 -5142 2417 -5102
rect -2575 -5482 2417 -5442
rect -2575 -10394 -2044 -5482
rect 1886 -10394 2417 -5482
rect -2575 -10434 2417 -10394
<< mimcap2contact >>
rect -2044 5482 1886 10394
rect -2044 190 1886 5102
rect -2044 -5102 1886 -190
rect -2044 -10394 1886 -5482
<< metal5 >>
rect -239 10418 81 10584
rect 2377 10493 2697 10584
rect -2068 10394 1910 10418
rect -2068 5482 -2044 10394
rect 1886 5482 1910 10394
rect -2068 5458 1910 5482
rect -239 5126 81 5458
rect 2377 5383 2419 10493
rect 2655 5383 2697 10493
rect 2377 5201 2697 5383
rect -2068 5102 1910 5126
rect -2068 190 -2044 5102
rect 1886 190 1910 5102
rect -2068 166 1910 190
rect -239 -166 81 166
rect 2377 91 2419 5201
rect 2655 91 2697 5201
rect 2377 -91 2697 91
rect -2068 -190 1910 -166
rect -2068 -5102 -2044 -190
rect 1886 -5102 1910 -190
rect -2068 -5126 1910 -5102
rect -239 -5458 81 -5126
rect 2377 -5201 2419 -91
rect 2655 -5201 2697 -91
rect 2377 -5383 2697 -5201
rect -2068 -5482 1910 -5458
rect -2068 -10394 -2044 -5482
rect 1886 -10394 1910 -5482
rect -2068 -10418 1910 -10394
rect -239 -10584 81 -10418
rect 2377 -10493 2419 -5383
rect 2655 -10493 2697 -5383
rect 2377 -10584 2697 -10493
<< properties >>
string FIXED_BBOX -2675 5342 2517 10534
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.962 l 24.962 val 1.265k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
