* NGSPICE file created from buffer.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_CL66SD a_1003_n100# a_803_n188# a_n2035_n188# a_n2711_n274#
+ a_n29_n100# a_487_n100# a_1835_n188# a_2293_n100# a_n229_n188# a_n1835_n100# a_287_n188#
+ a_n1003_n188# a_2093_n188# a_n803_n100# a_1519_n100# a_n2093_n100# a_1261_n100#
+ a_1319_n188# a_n2293_n188# a_n1319_n100# a_1061_n188# a_n287_n100# a_n1061_n100#
+ a_n1519_n188# a_745_n100# a_n487_n188# a_n1261_n188# a_2551_n100# a_545_n188# a_2351_n188#
+ a_1777_n100# a_n2609_n100# a_n2351_n100# a_1577_n188# a_229_n100# a_n1577_n100#
+ a_n2551_n188# a_2035_n100# a_n545_n100# a_n1777_n188# a_29_n188# a_n745_n188#
X0 a_n287_n100# a_n487_n188# a_n545_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_n2351_n100# a_n2551_n188# a_n2609_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X2 a_1777_n100# a_1577_n188# a_1519_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_2293_n100# a_2093_n188# a_2035_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_1003_n100# a_803_n188# a_745_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X5 a_n1577_n100# a_n1777_n188# a_n1835_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X6 a_n2093_n100# a_n2293_n188# a_n2351_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X7 a_n803_n100# a_n1003_n188# a_n1061_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X8 a_745_n100# a_545_n188# a_487_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X9 a_n29_n100# a_n229_n188# a_n287_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X10 a_229_n100# a_29_n188# a_n29_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X11 a_1519_n100# a_1319_n188# a_1261_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X12 a_487_n100# a_287_n188# a_229_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X13 a_n1319_n100# a_n1519_n188# a_n1577_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X14 a_n545_n100# a_n745_n188# a_n803_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X15 a_n1835_n100# a_n2035_n188# a_n2093_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X16 a_1261_n100# a_1061_n188# a_1003_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X17 a_2035_n100# a_1835_n188# a_1777_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X18 a_n1061_n100# a_n1261_n188# a_n1319_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X19 a_2551_n100# a_2351_n188# a_2293_n100# a_n2711_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
C0 a_n1261_n188# a_29_n188# 0.00fF
C1 a_n803_n100# a_n1577_n100# 0.00fF
C2 a_n803_n100# a_229_n100# 0.00fF
C3 a_487_n100# a_1061_n188# 0.00fF
C4 a_2093_n188# a_1261_n100# 0.00fF
C5 a_2551_n100# a_1519_n100# 0.00fF
C6 a_1003_n100# a_229_n100# 0.00fF
C7 a_n487_n188# a_n29_n100# 0.00fF
C8 a_n803_n100# a_n229_n188# 0.00fF
C9 a_29_n188# a_n1061_n100# 0.00fF
C10 a_1577_n188# a_287_n188# 0.00fF
C11 a_n745_n188# a_n803_n100# 0.00fF
C12 a_n487_n188# a_n287_n100# 0.00fF
C13 a_1003_n100# a_n229_n188# 0.00fF
C14 a_487_n100# a_n487_n188# 0.00fF
C15 a_1261_n100# a_n29_n100# 0.00fF
C16 a_803_n188# a_29_n188# 0.00fF
C17 a_1003_n100# a_745_n100# 0.06fF
C18 a_n2035_n188# a_n2293_n188# 0.10fF
C19 a_2351_n188# a_2551_n100# 0.00fF
C20 a_n1577_n100# a_n2093_n100# 0.00fF
C21 a_487_n100# a_1261_n100# 0.00fF
C22 a_n1319_n100# a_n2351_n100# 0.00fF
C23 a_n287_n100# a_n29_n100# 0.06fF
C24 a_487_n100# a_n29_n100# 0.00fF
C25 a_n2093_n100# a_n2551_n188# 0.00fF
C26 a_1777_n100# a_1319_n188# 0.00fF
C27 a_1319_n188# a_2035_n100# 0.00fF
C28 a_487_n100# a_n287_n100# 0.00fF
C29 a_n1319_n100# a_n545_n100# 0.00fF
C30 a_n487_n188# a_n1003_n188# 0.00fF
C31 a_1835_n188# a_545_n188# 0.00fF
C32 a_n1777_n188# a_n1003_n188# 0.00fF
C33 a_1319_n188# a_1519_n100# 0.00fF
C34 a_n803_n100# a_29_n188# 0.00fF
C35 a_545_n188# a_1577_n188# 0.00fF
C36 a_1003_n100# a_29_n188# 0.00fF
C37 a_n2609_n100# a_n1519_n188# 0.00fF
C38 a_n2035_n188# a_n2351_n100# 0.00fF
C39 a_n2293_n188# a_n2351_n100# 0.00fF
C40 a_n1003_n188# a_n29_n100# 0.00fF
C41 a_n1835_n100# a_n1777_n188# 0.00fF
C42 a_545_n188# a_287_n188# 0.10fF
C43 a_n1577_n100# a_n1319_n100# 0.06fF
C44 a_n287_n100# a_n1003_n188# 0.00fF
C45 a_803_n188# a_1319_n188# 0.00fF
C46 a_2351_n188# a_1319_n188# 0.00fF
C47 a_n1319_n100# a_n2551_n188# 0.00fF
C48 a_287_n188# a_n545_n100# 0.00fF
C49 a_2035_n100# a_2293_n100# 0.06fF
C50 a_1777_n100# a_2293_n100# 0.00fF
C51 a_n1319_n100# a_n229_n188# 0.00fF
C52 a_n745_n188# a_n1319_n100# 0.00fF
C53 a_1519_n100# a_2293_n100# 0.00fF
C54 a_1835_n188# a_745_n100# 0.00fF
C55 a_287_n188# a_229_n100# 0.00fF
C56 a_n2035_n188# a_n1577_n100# 0.00fF
C57 a_n1577_n100# a_n2293_n188# 0.00fF
C58 a_1003_n100# a_1319_n188# 0.00fF
C59 a_1577_n188# a_745_n100# 0.00fF
C60 a_n2035_n188# a_n2551_n188# 0.00fF
C61 a_n2551_n188# a_n2293_n188# 0.10fF
C62 a_287_n188# a_n229_n188# 0.00fF
C63 a_2351_n188# a_2293_n100# 0.00fF
C64 a_n745_n188# a_287_n188# 0.00fF
C65 a_n2035_n188# a_n745_n188# 0.00fF
C66 a_745_n100# a_287_n188# 0.00fF
C67 a_n1835_n100# a_n1003_n188# 0.00fF
C68 a_1777_n100# a_1061_n188# 0.00fF
C69 a_1061_n188# a_2035_n100# 0.00fF
C70 a_545_n188# a_n545_n100# 0.00fF
C71 a_1061_n188# a_1519_n100# 0.00fF
C72 a_n2093_n100# a_n2609_n100# 0.00fF
C73 a_2093_n188# a_2035_n100# 0.00fF
C74 a_1777_n100# a_2093_n188# 0.00fF
C75 a_2551_n100# a_1835_n188# 0.00fF
C76 a_n1577_n100# a_n2351_n100# 0.00fF
C77 a_n1261_n188# a_n487_n188# 0.00fF
C78 a_1777_n100# a_1261_n100# 0.00fF
C79 a_2035_n100# a_1261_n100# 0.00fF
C80 a_545_n188# a_229_n100# 0.00fF
C81 a_n1261_n188# a_n1777_n188# 0.00fF
C82 a_2551_n100# a_1577_n188# 0.00fF
C83 a_n2551_n188# a_n2351_n100# 0.00fF
C84 a_1003_n100# a_2293_n100# 0.00fF
C85 a_2093_n188# a_1519_n100# 0.00fF
C86 a_n487_n188# a_n1519_n188# 0.00fF
C87 a_803_n188# a_1061_n188# 0.10fF
C88 a_n1777_n188# a_n1519_n188# 0.10fF
C89 a_29_n188# a_287_n188# 0.10fF
C90 a_2351_n188# a_1061_n188# 0.00fF
C91 a_n545_n100# a_229_n100# 0.00fF
C92 a_n1577_n100# a_n545_n100# 0.00fF
C93 a_1261_n100# a_1519_n100# 0.06fF
C94 a_n487_n188# a_n1061_n100# 0.00fF
C95 a_545_n188# a_n229_n188# 0.00fF
C96 a_n745_n188# a_545_n188# 0.00fF
C97 a_n1777_n188# a_n1061_n100# 0.00fF
C98 a_487_n100# a_1777_n100# 0.00fF
C99 a_n1261_n188# a_n29_n100# 0.00fF
C100 a_545_n188# a_745_n100# 0.00fF
C101 a_803_n188# a_n487_n188# 0.00fF
C102 a_n545_n100# a_n229_n188# 0.00fF
C103 a_n1261_n188# a_n287_n100# 0.00fF
C104 a_n745_n188# a_n545_n100# 0.00fF
C105 a_803_n188# a_2093_n188# 0.00fF
C106 a_2351_n188# a_2093_n188# 0.10fF
C107 a_745_n100# a_n545_n100# 0.00fF
C108 a_487_n100# a_1519_n100# 0.00fF
C109 a_n1319_n100# a_n2609_n100# 0.00fF
C110 a_n287_n100# a_n1519_n188# 0.00fF
C111 a_n1061_n100# a_n29_n100# 0.00fF
C112 a_803_n188# a_1261_n100# 0.00fF
C113 a_2351_n188# a_1261_n100# 0.00fF
C114 a_n287_n100# a_n1061_n100# 0.00fF
C115 a_803_n188# a_n29_n100# 0.00fF
C116 a_1319_n188# a_1835_n188# 0.00fF
C117 a_n1577_n100# a_n2551_n188# 0.00fF
C118 a_1003_n100# a_1061_n188# 0.00fF
C119 a_n229_n188# a_229_n100# 0.00fF
C120 a_803_n188# a_n287_n100# 0.00fF
C121 a_n745_n188# a_n1577_n100# 0.00fF
C122 a_n745_n188# a_229_n100# 0.00fF
C123 a_803_n188# a_487_n100# 0.00fF
C124 a_1319_n188# a_1577_n188# 0.10fF
C125 a_745_n100# a_229_n100# 0.00fF
C126 a_29_n188# a_545_n188# 0.00fF
C127 a_n803_n100# a_n487_n188# 0.00fF
C128 a_n803_n100# a_n1777_n188# 0.00fF
C129 a_n1261_n188# a_n1003_n188# 0.10fF
C130 a_1319_n188# a_287_n188# 0.00fF
C131 a_1003_n100# a_2093_n188# 0.00fF
C132 a_n745_n188# a_n229_n188# 0.00fF
C133 a_n1003_n188# a_n1519_n188# 0.00fF
C134 a_29_n188# a_n545_n100# 0.00fF
C135 a_n2035_n188# a_n2609_n100# 0.00fF
C136 a_745_n100# a_n229_n188# 0.00fF
C137 a_n2293_n188# a_n2609_n100# 0.00fF
C138 a_1003_n100# a_1261_n100# 0.06fF
C139 a_n1061_n100# a_n1003_n188# 0.00fF
C140 a_n803_n100# a_n29_n100# 0.00fF
C141 a_n1261_n188# a_n1835_n100# 0.00fF
C142 a_1003_n100# a_n29_n100# 0.00fF
C143 a_n803_n100# a_n287_n100# 0.00fF
C144 a_n1835_n100# a_n1519_n188# 0.00fF
C145 a_487_n100# a_n803_n100# 0.00fF
C146 a_1835_n188# a_2293_n100# 0.00fF
C147 a_1003_n100# a_n287_n100# 0.00fF
C148 a_n2093_n100# a_n1777_n188# 0.00fF
C149 a_n1835_n100# a_n1061_n100# 0.00fF
C150 a_487_n100# a_1003_n100# 0.00fF
C151 a_29_n188# a_229_n100# 0.00fF
C152 a_1577_n188# a_2293_n100# 0.00fF
C153 a_29_n188# a_n229_n188# 0.10fF
C154 a_n745_n188# a_29_n188# 0.00fF
C155 a_n2609_n100# a_n2351_n100# 0.06fF
C156 a_1319_n188# a_545_n188# 0.00fF
C157 a_29_n188# a_745_n100# 0.00fF
C158 a_n803_n100# a_n1003_n188# 0.00fF
C159 a_n487_n188# a_n1319_n100# 0.00fF
C160 a_1835_n188# a_1061_n188# 0.00fF
C161 a_n1777_n188# a_n1319_n100# 0.00fF
C162 a_n1835_n100# a_n803_n100# 0.00fF
C163 a_1061_n188# a_1577_n188# 0.00fF
C164 a_1777_n100# a_2035_n100# 0.06fF
C165 a_1319_n188# a_229_n100# 0.00fF
C166 a_1835_n188# a_2093_n188# 0.10fF
C167 a_n2093_n100# a_n1003_n188# 0.00fF
C168 a_n1319_n100# a_n29_n100# 0.00fF
C169 a_1061_n188# a_287_n188# 0.00fF
C170 a_n1577_n100# a_n2609_n100# 0.00fF
C171 a_1777_n100# a_1519_n100# 0.06fF
C172 a_2035_n100# a_1519_n100# 0.00fF
C173 a_n287_n100# a_n1319_n100# 0.00fF
C174 a_1835_n188# a_1261_n100# 0.00fF
C175 a_2093_n188# a_1577_n188# 0.00fF
C176 a_n2551_n188# a_n2609_n100# 0.00fF
C177 a_n1835_n100# a_n2093_n100# 0.06fF
C178 a_n487_n188# a_287_n188# 0.00fF
C179 a_1261_n100# a_1577_n188# 0.00fF
C180 a_1319_n188# a_745_n100# 0.00fF
C181 a_n2035_n188# a_n1777_n188# 0.10fF
C182 a_n1261_n188# a_n1519_n188# 0.10fF
C183 a_n1777_n188# a_n2293_n188# 0.00fF
C184 a_1261_n100# a_287_n188# 0.00fF
C185 a_803_n188# a_1777_n100# 0.00fF
C186 a_803_n188# a_2035_n100# 0.00fF
C187 a_n1261_n188# a_n1061_n100# 0.00fF
C188 a_2351_n188# a_2035_n100# 0.00fF
C189 a_2351_n188# a_1777_n100# 0.00fF
C190 a_487_n100# a_1577_n188# 0.00fF
C191 a_n1061_n100# a_n1519_n188# 0.00fF
C192 a_287_n188# a_n29_n100# 0.00fF
C193 a_803_n188# a_1519_n100# 0.00fF
C194 a_n1319_n100# a_n1003_n188# 0.00fF
C195 a_n287_n100# a_287_n188# 0.00fF
C196 a_2351_n188# a_1519_n100# 0.00fF
C197 a_487_n100# a_287_n188# 0.00fF
C198 a_1061_n188# a_545_n188# 0.00fF
C199 a_1319_n188# a_29_n188# 0.00fF
C200 a_n1835_n100# a_n1319_n100# 0.00fF
C201 a_2551_n100# a_1319_n188# 0.00fF
C202 a_n1777_n188# a_n2351_n100# 0.00fF
C203 a_n487_n188# a_545_n188# 0.00fF
C204 a_1003_n100# a_2035_n100# 0.00fF
C205 a_1003_n100# a_1777_n100# 0.00fF
C206 a_n1261_n188# a_n803_n100# 0.00fF
C207 a_n487_n188# a_n545_n100# 0.00fF
C208 a_1261_n100# a_545_n188# 0.00fF
C209 a_287_n188# a_n1003_n188# 0.00fF
C210 a_n1777_n188# a_n545_n100# 0.00fF
C211 a_n2035_n188# a_n1003_n188# 0.00fF
C212 a_n803_n100# a_n1519_n188# 0.00fF
C213 a_n2293_n188# a_n1003_n188# 0.00fF
C214 a_1003_n100# a_1519_n100# 0.00fF
C215 a_545_n188# a_n29_n100# 0.00fF
C216 a_1061_n188# a_229_n100# 0.00fF
C217 a_n803_n100# a_n1061_n100# 0.06fF
C218 a_n287_n100# a_545_n188# 0.00fF
C219 a_487_n100# a_545_n188# 0.00fF
C220 a_n545_n100# a_n29_n100# 0.00fF
C221 a_n2035_n188# a_n1835_n100# 0.00fF
C222 a_n1835_n100# a_n2293_n188# 0.00fF
C223 a_1061_n188# a_n229_n188# 0.00fF
C224 a_n487_n188# a_229_n100# 0.00fF
C225 a_n1577_n100# a_n487_n188# 0.00fF
C226 a_n287_n100# a_n545_n100# 0.06fF
C227 a_n1577_n100# a_n1777_n188# 0.00fF
C228 a_n1261_n188# a_n2093_n100# 0.00fF
C229 a_803_n188# a_1003_n100# 0.00fF
C230 a_2551_n100# a_2293_n100# 0.06fF
C231 a_487_n100# a_n545_n100# 0.00fF
C232 a_1061_n188# a_745_n100# 0.00fF
C233 a_n2093_n100# a_n1519_n188# 0.00fF
C234 a_n1777_n188# a_n2551_n188# 0.00fF
C235 a_1261_n100# a_229_n100# 0.00fF
C236 a_n487_n188# a_n229_n188# 0.10fF
C237 a_n745_n188# a_n487_n188# 0.10fF
C238 a_n745_n188# a_n1777_n188# 0.00fF
C239 a_n2093_n100# a_n1061_n100# 0.00fF
C240 a_n487_n188# a_745_n100# 0.00fF
C241 a_229_n100# a_n29_n100# 0.06fF
C242 a_n1577_n100# a_n287_n100# 0.00fF
C243 a_n287_n100# a_229_n100# 0.00fF
C244 a_487_n100# a_229_n100# 0.06fF
C245 a_1261_n100# a_745_n100# 0.00fF
C246 a_n229_n188# a_n29_n100# 0.00fF
C247 a_n745_n188# a_n29_n100# 0.00fF
C248 a_n545_n100# a_n1003_n188# 0.00fF
C249 a_n1835_n100# a_n2351_n100# 0.00fF
C250 a_745_n100# a_n29_n100# 0.00fF
C251 a_n287_n100# a_n229_n188# 0.00fF
C252 a_29_n188# a_1061_n188# 0.00fF
C253 a_n745_n188# a_n287_n100# 0.00fF
C254 a_487_n100# a_n229_n188# 0.00fF
C255 a_n745_n188# a_487_n100# 0.00fF
C256 a_n1261_n188# a_n1319_n100# 0.00fF
C257 a_n287_n100# a_745_n100# 0.00fF
C258 a_487_n100# a_745_n100# 0.06fF
C259 a_1777_n100# a_1835_n188# 0.00fF
C260 a_1835_n188# a_2035_n100# 0.00fF
C261 a_n1319_n100# a_n1519_n188# 0.00fF
C262 a_n1835_n100# a_n545_n100# 0.00fF
C263 a_1319_n188# a_2293_n100# 0.00fF
C264 a_n487_n188# a_29_n188# 0.00fF
C265 a_1777_n100# a_1577_n188# 0.00fF
C266 a_2035_n100# a_1577_n188# 0.00fF
C267 a_n1319_n100# a_n1061_n100# 0.06fF
C268 a_n803_n100# a_n2093_n100# 0.00fF
C269 a_n1003_n188# a_229_n100# 0.00fF
C270 a_n1577_n100# a_n1003_n188# 0.00fF
C271 a_2551_n100# a_2093_n188# 0.00fF
C272 a_1835_n188# a_1519_n100# 0.00fF
C273 a_29_n188# a_1261_n100# 0.00fF
C274 a_2551_n100# a_1261_n100# 0.00fF
C275 a_1519_n100# a_1577_n188# 0.00fF
C276 a_n229_n188# a_n1003_n188# 0.00fF
C277 a_29_n188# a_n29_n100# 0.00fF
C278 a_n745_n188# a_n1003_n188# 0.10fF
C279 a_n1835_n100# a_n1577_n100# 0.06fF
C280 a_n2035_n188# a_n1261_n188# 0.00fF
C281 a_n1261_n188# a_n2293_n188# 0.00fF
C282 a_29_n188# a_n287_n100# 0.00fF
C283 a_1519_n100# a_287_n188# 0.00fF
C284 a_487_n100# a_29_n188# 0.00fF
C285 a_803_n188# a_1835_n188# 0.00fF
C286 a_n1835_n100# a_n2551_n188# 0.00fF
C287 a_2351_n188# a_1835_n188# 0.00fF
C288 a_n2035_n188# a_n1519_n188# 0.00fF
C289 a_n2293_n188# a_n1519_n188# 0.00fF
C290 a_n1835_n100# a_n745_n188# 0.00fF
C291 a_803_n188# a_1577_n188# 0.00fF
C292 a_1319_n188# a_1061_n188# 0.10fF
C293 a_n2035_n188# a_n1061_n100# 0.00fF
C294 a_2351_n188# a_1577_n188# 0.00fF
C295 a_n2293_n188# a_n1061_n100# 0.00fF
C296 a_n803_n100# a_n1319_n100# 0.00fF
C297 a_803_n188# a_287_n188# 0.00fF
C298 a_1319_n188# a_2093_n188# 0.00fF
C299 a_29_n188# a_n1003_n188# 0.00fF
C300 a_n1777_n188# a_n2609_n100# 0.00fF
C301 a_1777_n100# a_545_n188# 0.00fF
C302 a_n1261_n188# a_n2351_n100# 0.00fF
C303 a_1319_n188# a_1261_n100# 0.00fF
C304 a_1003_n100# a_1835_n188# 0.00fF
C305 a_n2351_n100# a_n1519_n188# 0.00fF
C306 a_545_n188# a_1519_n100# 0.00fF
C307 a_n2093_n100# a_n1319_n100# 0.00fF
C308 a_1003_n100# a_1577_n188# 0.00fF
C309 a_n1061_n100# a_n2351_n100# 0.00fF
C310 a_n803_n100# a_287_n188# 0.00fF
C311 a_n1261_n188# a_n545_n100# 0.00fF
C312 a_1061_n188# a_2293_n100# 0.00fF
C313 a_n2035_n188# a_n803_n100# 0.00fF
C314 a_487_n100# a_1319_n188# 0.00fF
C315 a_1003_n100# a_287_n188# 0.00fF
C316 a_n545_n100# a_n1519_n188# 0.00fF
C317 a_803_n188# a_545_n188# 0.10fF
C318 a_n545_n100# a_n1061_n100# 0.00fF
C319 a_2093_n188# a_2293_n100# 0.00fF
C320 a_n1261_n188# a_n1577_n100# 0.00fF
C321 a_1261_n100# a_2293_n100# 0.00fF
C322 a_1519_n100# a_229_n100# 0.00fF
C323 a_n2035_n188# a_n2093_n100# 0.00fF
C324 a_n1577_n100# a_n1519_n188# 0.00fF
C325 a_n2093_n100# a_n2293_n188# 0.00fF
C326 a_n1261_n188# a_n2551_n188# 0.00fF
C327 a_2035_n100# a_745_n100# 0.00fF
C328 a_1777_n100# a_745_n100# 0.00fF
C329 a_n1261_n188# a_n229_n188# 0.00fF
C330 a_n1261_n188# a_n745_n188# 0.00fF
C331 a_n2551_n188# a_n1519_n188# 0.00fF
C332 a_n1577_n100# a_n1061_n100# 0.00fF
C333 a_n1061_n100# a_229_n100# 0.00fF
C334 a_n229_n188# a_n1519_n188# 0.00fF
C335 a_n745_n188# a_n1519_n188# 0.00fF
C336 a_1519_n100# a_745_n100# 0.00fF
C337 a_803_n188# a_229_n100# 0.00fF
C338 a_1003_n100# a_545_n188# 0.00fF
C339 a_n229_n188# a_n1061_n100# 0.00fF
C340 a_n1835_n100# a_n2609_n100# 0.00fF
C341 a_n745_n188# a_n1061_n100# 0.00fF
C342 a_n803_n100# a_n545_n100# 0.06fF
C343 a_2093_n188# a_1061_n188# 0.00fF
C344 a_803_n188# a_n229_n188# 0.00fF
C345 a_803_n188# a_745_n100# 0.00fF
C346 a_1061_n188# a_1261_n100# 0.00fF
C347 a_n2093_n100# a_n2351_n100# 0.06fF
C348 a_n2035_n188# a_n1319_n100# 0.00fF
C349 a_n1319_n100# a_n2293_n188# 0.00fF
C350 a_2551_n100# a_2035_n100# 0.00fF
C351 a_2551_n100# a_1777_n100# 0.00fF
C352 a_n487_n188# a_n1777_n188# 0.00fF
C353 a_1835_n188# a_1577_n188# 0.10fF
C354 a_1061_n188# a_n29_n100# 0.00fF
C355 a_2551_n100# a_n2711_n274# 0.11fF
C356 a_2293_n100# a_n2711_n274# 0.05fF
C357 a_2035_n100# a_n2711_n274# 0.05fF
C358 a_1777_n100# a_n2711_n274# 0.04fF
C359 a_1519_n100# a_n2711_n274# 0.04fF
C360 a_1261_n100# a_n2711_n274# 0.04fF
C361 a_1003_n100# a_n2711_n274# 0.04fF
C362 a_745_n100# a_n2711_n274# 0.04fF
C363 a_487_n100# a_n2711_n274# 0.04fF
C364 a_229_n100# a_n2711_n274# 0.04fF
C365 a_n29_n100# a_n2711_n274# 0.04fF
C366 a_n287_n100# a_n2711_n274# 0.04fF
C367 a_n545_n100# a_n2711_n274# 0.04fF
C368 a_n803_n100# a_n2711_n274# 0.04fF
C369 a_n1061_n100# a_n2711_n274# 0.04fF
C370 a_n1319_n100# a_n2711_n274# 0.04fF
C371 a_n1577_n100# a_n2711_n274# 0.04fF
C372 a_n1835_n100# a_n2711_n274# 0.04fF
C373 a_n2093_n100# a_n2711_n274# 0.05fF
C374 a_n2351_n100# a_n2711_n274# 0.05fF
C375 a_n2609_n100# a_n2711_n274# 0.13fF
C376 a_2351_n188# a_n2711_n274# 0.63fF
C377 a_2093_n188# a_n2711_n274# 0.55fF
C378 a_1835_n188# a_n2711_n274# 0.55fF
C379 a_1577_n188# a_n2711_n274# 0.55fF
C380 a_1319_n188# a_n2711_n274# 0.54fF
C381 a_1061_n188# a_n2711_n274# 0.54fF
C382 a_803_n188# a_n2711_n274# 0.54fF
C383 a_545_n188# a_n2711_n274# 0.54fF
C384 a_287_n188# a_n2711_n274# 0.54fF
C385 a_29_n188# a_n2711_n274# 0.54fF
C386 a_n229_n188# a_n2711_n274# 0.54fF
C387 a_n487_n188# a_n2711_n274# 0.54fF
C388 a_n745_n188# a_n2711_n274# 0.54fF
C389 a_n1003_n188# a_n2711_n274# 0.54fF
C390 a_n1261_n188# a_n2711_n274# 0.54fF
C391 a_n1519_n188# a_n2711_n274# 0.54fF
C392 a_n1777_n188# a_n2711_n274# 0.55fF
C393 a_n2035_n188# a_n2711_n274# 0.55fF
C394 a_n2293_n188# a_n2711_n274# 0.55fF
C395 a_n2551_n188# a_n2711_n274# 0.63fF
.ends

.subckt sky130_fd_pr__pfet_01v8_BLSBYX w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
C0 a_n158_n100# w_n296_n319# 0.16fF
C1 a_100_n100# w_n296_n319# 0.07fF
C2 w_n296_n319# a_n100_n197# 0.29fF
C3 a_n158_n100# a_100_n100# 0.06fF
C4 a_100_n100# a_n100_n197# 0.00fF
C5 a_n158_n100# a_n100_n197# 0.00fF
C6 a_100_n100# VSUBS 0.06fF
C7 a_n158_n100# VSUBS 0.03fF
C8 a_n100_n197# VSUBS 0.36fF
C9 w_n296_n319# VSUBS 1.66fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8L4H97 a_158_n197# a_n416_n100# w_n812_n319# a_n358_n197#
+ a_358_n100# a_416_n197# a_n100_n197# a_100_n100# a_n674_n100# a_n158_n100# a_n616_n197#
+ a_616_n100# VSUBS
X0 a_n158_n100# a_n358_n197# a_n416_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X2 a_616_n100# a_416_n197# a_358_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_358_n100# a_158_n197# a_100_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4 a_n416_n100# a_n616_n197# a_n674_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
C0 a_416_n197# a_n616_n197# 0.00fF
C1 a_616_n100# a_n158_n100# 0.00fF
C2 a_100_n100# a_n674_n100# 0.00fF
C3 a_616_n100# a_358_n100# 0.03fF
C4 a_n416_n100# a_n158_n100# 0.03fF
C5 a_100_n100# a_416_n197# 0.00fF
C6 a_n416_n100# a_358_n100# 0.00fF
C7 a_n158_n100# a_358_n100# 0.01fF
C8 a_n100_n197# a_158_n197# 0.11fF
C9 a_n358_n197# a_158_n197# 0.00fF
C10 a_n616_n197# a_158_n197# 0.00fF
C11 a_100_n100# a_158_n197# 0.00fF
C12 a_n416_n100# a_n674_n100# 0.03fF
C13 a_416_n197# a_616_n100# 0.00fF
C14 a_n100_n197# w_n812_n319# 0.36fF
C15 a_n358_n197# w_n812_n319# 0.36fF
C16 a_416_n197# a_n416_n100# 0.00fF
C17 w_n812_n319# a_n616_n197# 0.39fF
C18 a_n158_n100# a_n674_n100# 0.01fF
C19 a_n674_n100# a_358_n100# 0.00fF
C20 a_416_n197# a_n158_n100# 0.00fF
C21 a_416_n197# a_358_n100# 0.00fF
C22 a_100_n100# w_n812_n319# 0.05fF
C23 a_616_n100# a_158_n197# 0.00fF
C24 a_n416_n100# a_158_n197# 0.00fF
C25 a_158_n197# a_n158_n100# 0.00fF
C26 a_416_n197# a_n674_n100# 0.00fF
C27 a_158_n197# a_358_n100# 0.00fF
C28 a_n358_n197# a_n100_n197# 0.11fF
C29 a_616_n100# w_n812_n319# 0.07fF
C30 a_n100_n197# a_n616_n197# 0.00fF
C31 a_n358_n197# a_n616_n197# 0.11fF
C32 a_n416_n100# w_n812_n319# 0.05fF
C33 a_100_n100# a_n100_n197# 0.00fF
C34 a_100_n100# a_n358_n197# 0.00fF
C35 w_n812_n319# a_n158_n100# 0.05fF
C36 a_100_n100# a_n616_n197# 0.00fF
C37 w_n812_n319# a_358_n100# 0.05fF
C38 a_158_n197# a_n674_n100# 0.00fF
C39 a_416_n197# a_158_n197# 0.11fF
C40 a_616_n100# a_n100_n197# 0.00fF
C41 a_n358_n197# a_616_n100# 0.00fF
C42 w_n812_n319# a_n674_n100# 0.09fF
C43 a_n416_n100# a_n358_n197# 0.00fF
C44 a_616_n100# a_n616_n197# 0.00fF
C45 a_n416_n100# a_n100_n197# 0.00fF
C46 a_416_n197# w_n812_n319# 0.39fF
C47 a_n416_n100# a_n616_n197# 0.00fF
C48 a_n100_n197# a_n158_n100# 0.00fF
C49 a_n358_n197# a_n158_n100# 0.00fF
C50 a_100_n100# a_616_n100# 0.01fF
C51 a_n100_n197# a_358_n100# 0.00fF
C52 a_n358_n197# a_358_n100# 0.00fF
C53 a_n616_n197# a_n158_n100# 0.00fF
C54 a_100_n100# a_n416_n100# 0.01fF
C55 a_n616_n197# a_358_n100# 0.00fF
C56 a_100_n100# a_n158_n100# 0.03fF
C57 a_100_n100# a_358_n100# 0.03fF
C58 w_n812_n319# a_158_n197# 0.36fF
C59 a_n100_n197# a_n674_n100# 0.00fF
C60 a_n358_n197# a_n674_n100# 0.00fF
C61 a_n616_n197# a_n674_n100# 0.00fF
C62 a_416_n197# a_n100_n197# 0.00fF
C63 a_416_n197# a_n358_n197# 0.00fF
C64 a_n416_n100# a_616_n100# 0.00fF
C65 a_616_n100# VSUBS 0.02fF
C66 a_358_n100# VSUBS 0.01fF
C67 a_100_n100# VSUBS 0.01fF
C68 a_n158_n100# VSUBS 0.01fF
C69 a_n416_n100# VSUBS 0.01fF
C70 a_n674_n100# VSUBS 0.02fF
C71 a_416_n197# VSUBS 0.27fF
C72 a_158_n197# VSUBS 0.22fF
C73 a_n100_n197# VSUBS 0.22fF
C74 a_n358_n197# VSUBS 0.22fF
C75 a_n616_n197# VSUBS 0.27fF
C76 w_n812_n319# VSUBS 4.34fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8C4HA7 a_158_n197# a_n416_n100# w_n812_n319# a_n358_n197#
+ a_358_n100# a_416_n197# a_n100_n197# a_100_n100# a_n674_n100# a_n158_n100# a_n616_n197#
+ a_616_n100# VSUBS
X0 a_n158_n100# a_n358_n197# a_n416_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X2 a_616_n100# a_416_n197# a_358_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_358_n100# a_158_n197# a_100_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4 a_n416_n100# a_n616_n197# a_n674_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
C0 a_616_n100# a_n358_n197# 0.00fF
C1 a_616_n100# a_n158_n100# 0.00fF
C2 a_616_n100# a_158_n197# 0.00fF
C3 a_n416_n100# a_100_n100# 0.01fF
C4 a_n100_n197# a_n674_n100# 0.00fF
C5 a_416_n197# a_n358_n197# 0.00fF
C6 a_416_n197# a_n158_n100# 0.00fF
C7 a_416_n197# a_158_n197# 0.11fF
C8 a_n616_n197# a_n358_n197# 0.11fF
C9 a_n616_n197# a_n158_n100# 0.00fF
C10 a_n100_n197# w_n812_n319# 0.36fF
C11 a_n616_n197# a_158_n197# 0.00fF
C12 a_n100_n197# a_n416_n100# 0.00fF
C13 a_n358_n197# a_n158_n100# 0.00fF
C14 a_n358_n197# a_158_n197# 0.00fF
C15 a_158_n197# a_n158_n100# 0.00fF
C16 a_616_n100# w_n812_n319# 0.07fF
C17 a_416_n197# a_n674_n100# 0.00fF
C18 a_616_n100# a_n416_n100# 0.00fF
C19 a_n616_n197# a_n674_n100# 0.00fF
C20 w_n812_n319# a_416_n197# 0.39fF
C21 w_n812_n319# a_n616_n197# 0.39fF
C22 a_416_n197# a_n416_n100# 0.00fF
C23 a_n358_n197# a_n674_n100# 0.00fF
C24 a_n674_n100# a_n158_n100# 0.01fF
C25 a_n674_n100# a_158_n197# 0.00fF
C26 a_n616_n197# a_n416_n100# 0.00fF
C27 w_n812_n319# a_n358_n197# 0.36fF
C28 w_n812_n319# a_n158_n100# 0.05fF
C29 w_n812_n319# a_158_n197# 0.36fF
C30 a_n416_n100# a_n358_n197# 0.00fF
C31 a_n416_n100# a_n158_n100# 0.03fF
C32 a_n416_n100# a_158_n197# 0.00fF
C33 a_358_n100# a_100_n100# 0.03fF
C34 w_n812_n319# a_n674_n100# 0.09fF
C35 a_n100_n197# a_358_n100# 0.00fF
C36 a_n416_n100# a_n674_n100# 0.03fF
C37 w_n812_n319# a_n416_n100# 0.05fF
C38 a_n100_n197# a_100_n100# 0.00fF
C39 a_616_n100# a_358_n100# 0.03fF
C40 a_358_n100# a_416_n197# 0.00fF
C41 a_616_n100# a_100_n100# 0.01fF
C42 a_358_n100# a_n616_n197# 0.00fF
C43 a_416_n197# a_100_n100# 0.00fF
C44 a_n616_n197# a_100_n100# 0.00fF
C45 a_358_n100# a_n358_n197# 0.00fF
C46 a_358_n100# a_n158_n100# 0.01fF
C47 a_358_n100# a_158_n197# 0.00fF
C48 a_n100_n197# a_616_n100# 0.00fF
C49 a_100_n100# a_n358_n197# 0.00fF
C50 a_100_n100# a_n158_n100# 0.03fF
C51 a_100_n100# a_158_n197# 0.00fF
C52 a_n100_n197# a_416_n197# 0.00fF
C53 a_n100_n197# a_n616_n197# 0.00fF
C54 a_n100_n197# a_n358_n197# 0.11fF
C55 a_n100_n197# a_n158_n100# 0.00fF
C56 a_n100_n197# a_158_n197# 0.11fF
C57 a_358_n100# a_n674_n100# 0.00fF
C58 a_616_n100# a_416_n197# 0.00fF
C59 a_358_n100# w_n812_n319# 0.05fF
C60 a_616_n100# a_n616_n197# 0.00fF
C61 a_100_n100# a_n674_n100# 0.00fF
C62 a_358_n100# a_n416_n100# 0.00fF
C63 w_n812_n319# a_100_n100# 0.05fF
C64 a_n616_n197# a_416_n197# 0.00fF
C65 a_616_n100# VSUBS 0.02fF
C66 a_358_n100# VSUBS 0.01fF
C67 a_100_n100# VSUBS 0.01fF
C68 a_n158_n100# VSUBS 0.01fF
C69 a_n416_n100# VSUBS 0.01fF
C70 a_n674_n100# VSUBS 0.02fF
C71 a_416_n197# VSUBS 0.27fF
C72 a_158_n197# VSUBS 0.22fF
C73 a_n100_n197# VSUBS 0.22fF
C74 a_n358_n197# VSUBS 0.22fF
C75 a_n616_n197# VSUBS 0.27fF
C76 w_n812_n319# VSUBS 4.34fF
.ends

.subckt sky130_fd_pr__nfet_01v8_GVTB53 a_n29_n100# a_n229_n188# a_n389_n274# a_n287_n100#
+ a_229_n100# a_29_n188#
X0 a_n29_n100# a_n229_n188# a_n287_n100# a_n389_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_229_n100# a_29_n188# a_n29_n100# a_n389_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
C0 a_29_n188# a_n29_n100# 0.00fF
C1 a_n229_n188# a_n287_n100# 0.00fF
C2 a_n229_n188# a_29_n188# 0.10fF
C3 a_29_n188# a_n287_n100# 0.00fF
C4 a_229_n100# a_n29_n100# 0.06fF
C5 a_229_n100# a_n229_n188# 0.00fF
C6 a_n229_n188# a_n29_n100# 0.00fF
C7 a_229_n100# a_n287_n100# 0.00fF
C8 a_n29_n100# a_n287_n100# 0.06fF
C9 a_229_n100# a_29_n188# 0.00fF
C10 a_229_n100# a_n389_n274# 0.13fF
C11 a_n29_n100# a_n389_n274# 0.08fF
C12 a_n287_n100# a_n389_n274# 0.15fF
C13 a_29_n188# a_n389_n274# 0.70fF
C14 a_n229_n188# a_n389_n274# 0.70fF
.ends

.subckt sky130_fd_pr__pfet_01v8_8LYGA7 a_158_n197# a_n416_n100# w_n812_n319# a_n358_n197#
+ a_358_n100# a_416_n197# a_n100_n197# a_100_n100# a_n674_n100# a_n158_n100# a_n616_n197#
+ a_616_n100# VSUBS
X0 a_n158_n100# a_n358_n197# a_n416_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X2 a_616_n100# a_416_n197# a_358_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_358_n100# a_158_n197# a_100_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4 a_n416_n100# a_n616_n197# a_n674_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
C0 a_416_n197# a_n358_n197# 0.00fF
C1 a_n416_n100# w_n812_n319# 0.04fF
C2 a_n616_n197# a_n100_n197# 0.00fF
C3 a_n100_n197# a_n158_n100# 0.00fF
C4 a_358_n100# a_n616_n197# 0.00fF
C5 a_358_n100# a_n158_n100# 0.01fF
C6 w_n812_n319# a_100_n100# 0.04fF
C7 w_n812_n319# a_n358_n197# 0.25fF
C8 a_n416_n100# a_100_n100# 0.01fF
C9 a_n416_n100# a_n358_n197# 0.00fF
C10 a_100_n100# a_n358_n197# 0.00fF
C11 a_416_n197# a_n674_n100# 0.00fF
C12 w_n812_n319# a_n674_n100# 0.12fF
C13 a_416_n197# a_n616_n197# 0.00fF
C14 a_416_n197# a_n158_n100# 0.00fF
C15 a_n416_n100# a_n674_n100# 0.03fF
C16 w_n812_n319# a_n616_n197# 0.30fF
C17 w_n812_n319# a_n158_n100# 0.04fF
C18 a_100_n100# a_n674_n100# 0.00fF
C19 a_n674_n100# a_n358_n197# 0.00fF
C20 a_n416_n100# a_n158_n100# 0.03fF
C21 a_n416_n100# a_n616_n197# 0.00fF
C22 a_158_n197# a_616_n100# 0.00fF
C23 a_100_n100# a_n616_n197# 0.00fF
C24 a_100_n100# a_n158_n100# 0.03fF
C25 a_n616_n197# a_n358_n197# 0.11fF
C26 a_n358_n197# a_n158_n100# 0.00fF
C27 a_616_n100# a_n100_n197# 0.00fF
C28 a_358_n100# a_616_n100# 0.03fF
C29 a_158_n197# a_n100_n197# 0.11fF
C30 a_358_n100# a_158_n197# 0.00fF
C31 a_358_n100# a_n100_n197# 0.00fF
C32 a_n674_n100# a_n158_n100# 0.01fF
C33 a_n616_n197# a_n674_n100# 0.00fF
C34 a_416_n197# a_616_n100# 0.00fF
C35 a_n616_n197# a_n158_n100# 0.00fF
C36 a_416_n197# a_158_n197# 0.11fF
C37 a_616_n100# w_n812_n319# 0.06fF
C38 a_158_n197# w_n812_n319# 0.25fF
C39 a_416_n197# a_n100_n197# 0.00fF
C40 a_358_n100# a_416_n197# 0.00fF
C41 a_n416_n100# a_616_n100# 0.00fF
C42 a_158_n197# a_n416_n100# 0.00fF
C43 a_616_n100# a_100_n100# 0.01fF
C44 a_616_n100# a_n358_n197# 0.00fF
C45 w_n812_n319# a_n100_n197# 0.25fF
C46 a_358_n100# w_n812_n319# 0.04fF
C47 a_158_n197# a_100_n100# 0.00fF
C48 a_158_n197# a_n358_n197# 0.00fF
C49 a_n416_n100# a_n100_n197# 0.00fF
C50 a_358_n100# a_n416_n100# 0.00fF
C51 a_100_n100# a_n100_n197# 0.00fF
C52 a_358_n100# a_100_n100# 0.03fF
C53 a_n100_n197# a_n358_n197# 0.11fF
C54 a_358_n100# a_n358_n197# 0.00fF
C55 a_158_n197# a_n674_n100# 0.00fF
C56 a_416_n197# w_n812_n319# 0.27fF
C57 a_616_n100# a_n616_n197# 0.00fF
C58 a_616_n100# a_n158_n100# 0.00fF
C59 a_n100_n197# a_n674_n100# 0.00fF
C60 a_358_n100# a_n674_n100# 0.00fF
C61 a_416_n197# a_n416_n100# 0.00fF
C62 a_158_n197# a_n616_n197# 0.00fF
C63 a_158_n197# a_n158_n100# 0.00fF
C64 a_416_n197# a_100_n100# 0.00fF
C65 a_616_n100# VSUBS 0.03fF
C66 a_358_n100# VSUBS 0.02fF
C67 a_100_n100# VSUBS 0.01fF
C68 a_n158_n100# VSUBS 0.01fF
C69 a_n416_n100# VSUBS 0.01fF
C70 a_n674_n100# VSUBS 0.01fF
C71 a_416_n197# VSUBS 0.30fF
C72 a_158_n197# VSUBS 0.24fF
C73 a_n100_n197# VSUBS 0.24fF
C74 a_n358_n197# VSUBS 0.24fF
C75 a_n616_n197# VSUBS 0.29fF
C76 w_n812_n319# VSUBS 4.13fF
.ends

.subckt buffer ib out in gnd vd
Xsky130_fd_pr__nfet_01v8_CL66SD_0 net2 out out gnd net2 net3 out net4 out net4 in
+ out out net4 net3 net2 net4 in out net4 out net4 net2 in net4 in out net3 in in
+ net4 net3 net4 in net4 net3 in net2 net3 in out in sky130_fd_pr__nfet_01v8_CL66SD
Xsky130_fd_pr__nfet_01v8_CL66SD_1 gnd net1 net1 gnd gnd gnd net1 out net1 out net1
+ net1 net1 out gnd gnd out net1 net1 net1 net1 net1 gnd net1 net1 net1 net1 gnd net1
+ net1 net1 gnd net1 net1 out gnd net1 gnd gnd net1 net1 net1 sky130_fd_pr__nfet_01v8_CL66SD
Xsky130_fd_pr__pfet_01v8_BLSBYX_0 vd net2 net2 vd gnd sky130_fd_pr__pfet_01v8_BLSBYX
Xsky130_fd_pr__pfet_01v8_8L4H97_0 net2 net1 vd net2 vd net2 net2 net1 vd vd net2 net1
+ gnd sky130_fd_pr__pfet_01v8_8L4H97
Xsky130_fd_pr__pfet_01v8_BLSBYX_1 vd net3 net3 vd gnd sky130_fd_pr__pfet_01v8_BLSBYX
Xsky130_fd_pr__pfet_01v8_8C4HA7_0 net3 out vd net3 vd net3 net3 out vd vd net3 out
+ gnd sky130_fd_pr__pfet_01v8_8C4HA7
Xsky130_fd_pr__nfet_01v8_GVTB53_0 gnd ib gnd ib net4 ib sky130_fd_pr__nfet_01v8_GVTB53
Xsky130_fd_pr__pfet_01v8_8LYGA7_0 net2 net1 vd net2 vd net2 net2 net1 vd vd net2 net1
+ gnd sky130_fd_pr__pfet_01v8_8LYGA7
Xsky130_fd_pr__pfet_01v8_8LYGA7_1 net3 out vd net3 vd net3 net3 out vd vd net3 out
+ gnd sky130_fd_pr__pfet_01v8_8LYGA7
X0 net2 out.t8 net4 gnd sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.29e+07u as=3.19e+12p ps=2.838e+07u w=0u l=0u
X1 net4 in.t2 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.548e+07u w=0u l=0u
X2 net4 in.t1 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X3 net2 out.t4 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X4 vd net2.t7 net1 vd sky130_fd_pr__pfet_01v8 ad=4.06e+12p pd=3.612e+07u as=1.74e+12p ps=1.548e+07u w=0u l=0u
X5 net4 out.t0 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X6 net3 in.t6 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X7 net3 in.t9 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X8 net4 out.t5 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X9 net4 out.t6 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X10 net2.t1 net2.t0 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X11 net1 net2.t9 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X12 net2 out.t2 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X13 net4 in.t0 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X14 gnd ib.t0 ib.t1 gnd sky130_fd_pr__nfet_01v8 ad=3.48e+12p pd=3.096e+07u as=0p ps=0u w=0u l=0u
X15 net4 ib.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X16 net3 in.t3 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X17 net4 out.t7 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X18 net4 in.t7 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X19 net2 out.t9 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X20 net4 in.t4 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X21 vd net2.t2 net1 vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X22 net1 net2.t6 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X23 net3 in.t5 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X24 net3 in.t8 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X25 net4 out.t3 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X26 net1 net2.t11 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X27 net2 out.t1 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X28 vd net2.t5 net1 vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X29 net1 net2.t3 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X30 net1 net2.t8 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X31 vd net2.t10 net1 vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
X32 net1 net2.t4 vd vd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=0u l=0u
R0 in.n1 in.n0 150.875
R1 in.n5 in.n4 150.49
R2 in.n3 in.n2 150.488
R3 in.n7 in.n6 141.16
R4 in.n0 in.t9 25.228
R5 in.n6 in.t7 24.105
R6 in.n0 in.t2 24.104
R7 in.n2 in.t4 24.103
R8 in.n4 in.t0 24.102
R9 in.n1 in.t5 24.102
R10 in.n5 in.t8 24.102
R11 in.n3 in.t6 24.102
R12 in.n7 in.t3 24.102
R13 in.n9 in.t1 24.1
R14 in.n14 in.n13 9.3
R15 in in.n14 5.261
R16 in.n8 in.n7 1.785
R17 in.n2 in.n1 1.103
R18 in.n4 in.n3 1.094
R19 in.n6 in.n5 0.41
R20 in.n14 in.n12 0.076
R21 in.n12 in.n8 0.014
R22 in.n12 in.n11 0.005
R23 in.n10 in.n9 0.005
R24 in.n11 in.n10 0.001
R25 out.t0 out.n7 175.091
R26 out.n0 out.t2 175.044
R27 out.n2 out.n1 150.491
R28 out.n4 out.n3 150.491
R29 out.n6 out.n5 141.106
R30 out out.t0 26.91
R31 out.n5 out.t1 24.103
R32 out.n6 out.t7 24.103
R33 out.n4 out.t5 24.103
R34 out.n2 out.t3 24.102
R35 out.n0 out.t6 24.102
R36 out.n1 out.t9 24.102
R37 out.n3 out.t4 24.102
R38 out.n7 out.t8 24.102
R39 out.n7 out.n6 1.085
R40 out.n3 out.n2 0.988
R41 out.n5 out.n4 0.913
R42 out.n1 out.n0 0.863
R43 net2.n4 net2.t6 40.035
R44 net2.n0 net2.t11 40.035
R45 net2.n8 net2.t0 39.528
R46 net2.n7 net2.t4 39.528
R47 net2.n6 net2.t5 39.528
R48 net2.n5 net2.t3 39.528
R49 net2.n4 net2.t2 39.528
R50 net2.n3 net2.t9 39.528
R51 net2.n2 net2.t10 39.528
R52 net2.n1 net2.t8 39.528
R53 net2.n0 net2.t7 39.528
R54 net2.n10 net2.t1 28.57
R55 net2.n8 net2.n7 1.982
R56 net2.n9 net2.n3 1.708
R57 net2 net2.n10 0.985
R58 net2.n5 net2.n4 0.507
R59 net2.n6 net2.n5 0.507
R60 net2.n7 net2.n6 0.507
R61 net2.n1 net2.n0 0.507
R62 net2.n2 net2.n1 0.507
R63 net2.n3 net2.n2 0.507
R64 net2.n10 net2.n9 0.335
R65 net2.n9 net2.n8 0.303
R66 vd.n53 vd.n52 379.482
R67 vd.n40 vd.n34 379.482
R68 vd.n54 vd.n53 297.411
R69 vd.n41 vd.n40 297.411
R70 vd.n19 vd.n16 131.387
R71 vd.n4 vd.n1 131.387
R72 vd.n24 vd.n21 131.011
R73 vd.n9 vd.n6 131.011
R74 vd.n29 vd.n24 54.211
R75 vd.n14 vd.n9 54.211
R76 vd.n29 vd.n19 53.835
R77 vd.n14 vd.n4 53.835
R78 vd.n57 vd.n14 8.271
R79 vd.n57 vd.n29 7.938
R80 vd.n57 vd.n56 4.028
R81 vd.n55 vd.n45 0.296
R82 vd vd.n57 0.28
R83 vd.n42 vd.n32 0.228
R84 vd.n56 vd.n55 0.18
R85 vd.n56 vd.n42 0.167
R86 vd.n19 vd.n18 0.161
R87 vd.n24 vd.n23 0.161
R88 vd.n4 vd.n3 0.161
R89 vd.n9 vd.n8 0.161
R90 vd.n23 vd.n22 0.139
R91 vd.n8 vd.n7 0.139
R92 vd.n18 vd.n17 0.139
R93 vd.n3 vd.n2 0.139
R94 vd.n42 vd.n41 0.017
R95 vd.n55 vd.n54 0.017
R96 vd.n16 vd.n15 0.015
R97 vd.n21 vd.n20 0.015
R98 vd.n1 vd.n0 0.015
R99 vd.n6 vd.n5 0.015
R100 vd.n52 vd.n51 0.013
R101 vd.n34 vd.n33 0.013
R102 vd.n26 vd.n25 0.013
R103 vd.n27 vd.n26 0.013
R104 vd.n11 vd.n10 0.013
R105 vd.n12 vd.n11 0.013
R106 vd.n53 vd.n50 0.003
R107 vd.n47 vd.n46 0.003
R108 vd.n36 vd.n35 0.003
R109 vd.n40 vd.n39 0.003
R110 vd.n50 vd.n49 0.003
R111 vd.n37 vd.n36 0.003
R112 vd.n48 vd.n47 0.003
R113 vd.n39 vd.n38 0.003
R114 vd.n49 vd.n48 0.002
R115 vd.n38 vd.n37 0.002
R116 vd.n29 vd.n28 0.002
R117 vd.n28 vd.n27 0.002
R118 vd.n14 vd.n13 0.002
R119 vd.n13 vd.n12 0.002
R120 vd.n32 vd.n31 0.001
R121 vd.n45 vd.n44 0.001
R122 vd.n44 vd.n43 0.001
R123 vd.n31 vd.n30 0.001
R124 ib.n0 ib.t2 24.837
R125 ib.n0 ib.t0 24.107
R126 ib.n1 ib.t1 17.747
R127 ib ib.n1 1.062
R128 ib.n1 ib.n0 0.387
C0 in net1 0.88fF
C1 net1 out 1.67fF
C2 in out 1.39fF
C3 net1 net4 0.18fF
C4 ib net1 0.04fF
C5 net3 net1 0.47fF
C6 in net4 2.12fF
C7 out net4 2.13fF
C8 ib in 0.06fF
C9 ib out 0.00fF
C10 vd net1 2.04fF
C11 net3 in 1.40fF
C12 net3 out 2.33fF
C13 in vd 0.81fF
C14 vd out 1.79fF
C15 ib net4 0.04fF
C16 net3 net4 2.19fF
C17 net3 ib 0.01fF
C18 net2 net1 2.18fF
C19 vd net4 0.09fF
C20 ib vd 0.02fF
C21 net3 vd 3.38fF
C22 net2 in 0.55fF
C23 net2 out 2.13fF
C24 net2 net4 1.85fF
C25 net3 net2 0.62fF
C26 net2 vd 4.36fF
C27 vd.n0 gnd 0.41fF $ **FLOATING
C28 vd.n1 gnd 0.07fF $ **FLOATING
C29 vd.n2 gnd 0.39fF $ **FLOATING
C30 vd.n3 gnd 0.04fF $ **FLOATING
C31 vd.n4 gnd 0.04fF $ **FLOATING
C32 vd.n5 gnd 0.41fF $ **FLOATING
C33 vd.n6 gnd 0.07fF $ **FLOATING
C34 vd.n7 gnd 0.39fF $ **FLOATING
C35 vd.n8 gnd 0.04fF $ **FLOATING
C36 vd.n9 gnd 0.04fF $ **FLOATING
C37 vd.n10 gnd 0.09fF $ **FLOATING
C38 vd.n11 gnd 0.09fF $ **FLOATING
C39 vd.n12 gnd 0.43fF $ **FLOATING
C40 vd.n13 gnd 0.02fF $ **FLOATING
C41 vd.n14 gnd 0.59fF $ **FLOATING
C42 vd.n15 gnd 0.41fF $ **FLOATING
C43 vd.n16 gnd 0.07fF $ **FLOATING
C44 vd.n17 gnd 0.39fF $ **FLOATING
C45 vd.n18 gnd 0.04fF $ **FLOATING
C46 vd.n19 gnd 0.04fF $ **FLOATING
C47 vd.n20 gnd 0.41fF $ **FLOATING
C48 vd.n21 gnd 0.07fF $ **FLOATING
C49 vd.n22 gnd 0.39fF $ **FLOATING
C50 vd.n23 gnd 0.04fF $ **FLOATING
C51 vd.n24 gnd 0.04fF $ **FLOATING
C52 vd.n25 gnd 0.09fF $ **FLOATING
C53 vd.n26 gnd 0.09fF $ **FLOATING
C54 vd.n27 gnd 0.43fF $ **FLOATING
C55 vd.n28 gnd 0.02fF $ **FLOATING
C56 vd.n29 gnd 0.62fF $ **FLOATING
C57 vd.n30 gnd 1.56fF $ **FLOATING
C58 vd.n31 gnd 0.04fF $ **FLOATING
C59 vd.n32 gnd 0.77fF $ **FLOATING
C60 vd.n33 gnd 1.56fF $ **FLOATING
C61 vd.n34 gnd 0.18fF $ **FLOATING
C62 vd.n35 gnd 0.15fF $ **FLOATING
C63 vd.n36 gnd 0.17fF $ **FLOATING
C64 vd.n37 gnd 1.21fF $ **FLOATING
C65 vd.n38 gnd 1.21fF $ **FLOATING
C66 vd.n39 gnd 0.17fF $ **FLOATING
C67 vd.n40 gnd 0.15fF $ **FLOATING
C68 vd.n41 gnd 0.09fF $ **FLOATING
C69 vd.n42 gnd 0.12fF $ **FLOATING
C70 vd.n43 gnd 1.56fF $ **FLOATING
C71 vd.n44 gnd 0.04fF $ **FLOATING
C72 vd.n45 gnd 0.41fF $ **FLOATING
C73 vd.n46 gnd 0.15fF $ **FLOATING
C74 vd.n47 gnd 0.17fF $ **FLOATING
C75 vd.n48 gnd 1.21fF $ **FLOATING
C76 vd.n49 gnd 1.21fF $ **FLOATING
C77 vd.n50 gnd 0.17fF $ **FLOATING
C78 vd.n51 gnd 1.56fF $ **FLOATING
C79 vd.n52 gnd 0.18fF $ **FLOATING
C80 vd.n53 gnd 0.15fF $ **FLOATING
C81 vd.n54 gnd 0.09fF $ **FLOATING
C82 vd.n55 gnd 0.42fF $ **FLOATING
C83 vd.n56 gnd 1.70fF $ **FLOATING
C84 vd.n57 gnd 15.86fF $ **FLOATING
C85 net2.t11 gnd 0.65fF
C86 net2.t7 gnd 0.65fF
C87 net2.n0 gnd 0.82fF $ **FLOATING
C88 net2.t8 gnd 0.65fF
C89 net2.n1 gnd 0.42fF $ **FLOATING
C90 net2.t10 gnd 0.65fF
C91 net2.n2 gnd 0.42fF $ **FLOATING
C92 net2.t9 gnd 0.65fF
C93 net2.n3 gnd 0.53fF $ **FLOATING
C94 net2.t0 gnd 0.65fF
C95 net2.t4 gnd 0.65fF
C96 net2.t5 gnd 0.65fF
C97 net2.t3 gnd 0.65fF
C98 net2.t2 gnd 0.65fF
C99 net2.t6 gnd 0.65fF
C100 net2.n4 gnd 0.82fF $ **FLOATING
C101 net2.n5 gnd 0.42fF $ **FLOATING
C102 net2.n6 gnd 0.42fF $ **FLOATING
C103 net2.n7 gnd 0.56fF $ **FLOATING
C104 net2.n8 gnd 0.53fF $ **FLOATING
C105 net2.n9 gnd 0.23fF $ **FLOATING
C106 net2.t1 gnd 0.03fF
C107 net2.n10 gnd 0.37fF $ **FLOATING
C108 out.t8 gnd 0.59fF
C109 out.t1 gnd 0.59fF
C110 out.t4 gnd 0.59fF
C111 out.t9 gnd 0.59fF
C112 out.t2 gnd 0.95fF
C113 out.t6 gnd 0.59fF
C114 out.n0 gnd 2.73fF $ **FLOATING
C115 out.n1 gnd 2.86fF $ **FLOATING
C116 out.t3 gnd 0.59fF
C117 out.n2 gnd 0.87fF $ **FLOATING
C118 out.n3 gnd 0.87fF $ **FLOATING
C119 out.t5 gnd 0.59fF
C120 out.n4 gnd 0.92fF $ **FLOATING
C121 out.n5 gnd 0.93fF $ **FLOATING
C122 out.t7 gnd 0.59fF
C123 out.n6 gnd 0.85fF $ **FLOATING
C124 out.n7 gnd 0.92fF $ **FLOATING
C125 out.t0 gnd 0.62fF
C126 in.t0 gnd 0.41fF
C127 in.t5 gnd 0.41fF
C128 in.t9 gnd 0.44fF
C129 in.t2 gnd 0.41fF
C130 in.n0 gnd 1.13fF $ **FLOATING
C131 in.n1 gnd 0.58fF $ **FLOATING
C132 in.t4 gnd 0.41fF
C133 in.n2 gnd 0.58fF $ **FLOATING
C134 in.t6 gnd 0.41fF
C135 in.n3 gnd 0.59fF $ **FLOATING
C136 in.n4 gnd 0.58fF $ **FLOATING
C137 in.t8 gnd 0.41fF
C138 in.n5 gnd 0.69fF $ **FLOATING
C139 in.t7 gnd 0.41fF
C140 in.n6 gnd 0.69fF $ **FLOATING
C141 in.t3 gnd 0.41fF
C142 in.n7 gnd 0.49fF $ **FLOATING
C143 in.n8 gnd 0.22fF $ **FLOATING
C144 in.t1 gnd 0.41fF
C145 in.n9 gnd 0.17fF $ **FLOATING
C146 in.n10 gnd 0.00fF $ **FLOATING
C147 in.n11 gnd 0.01fF $ **FLOATING
C148 in.n12 gnd 0.02fF $ **FLOATING
C149 in.n13 gnd 0.02fF $ **FLOATING
C150 in.n14 gnd 0.25fF $ **FLOATING
C151 net4 gnd 1.49fF
C152 ib gnd 1.87fF
C153 out gnd 13.46fF
C154 net3 gnd 3.38fF
C155 vd gnd 18.59fF
C156 net1 gnd 17.83fF
C157 net2 gnd 8.89fF
C158 in gnd 6.08fF
.ends

