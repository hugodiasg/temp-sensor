magic
tech sky130A
magscale 1 2
timestamp 1644769315
<< metal4 >>
rect -2519 7379 2519 7420
rect -2519 2581 2263 7379
rect 2499 2581 2519 7379
rect -2519 2540 2519 2581
rect -2519 2399 2519 2440
rect -2519 -2399 2263 2399
rect 2499 -2399 2519 2399
rect -2519 -2440 2519 -2399
rect -2519 -2581 2519 -2540
rect -2519 -7379 2263 -2581
rect 2499 -7379 2519 -2581
rect -2519 -7420 2519 -7379
<< via4 >>
rect 2263 2581 2499 7379
rect 2263 -2399 2499 2399
rect 2263 -7379 2499 -2581
<< mimcap2 >>
rect -2419 7280 2261 7320
rect -2419 2680 -1919 7280
rect 1761 2680 2261 7280
rect -2419 2640 2261 2680
rect -2419 2300 2261 2340
rect -2419 -2300 -1919 2300
rect 1761 -2300 2261 2300
rect -2419 -2340 2261 -2300
rect -2419 -2680 2261 -2640
rect -2419 -7280 -1919 -2680
rect 1761 -7280 2261 -2680
rect -2419 -7320 2261 -7280
<< mimcap2contact >>
rect -1919 2680 1761 7280
rect -1919 -2300 1761 2300
rect -1919 -7280 1761 -2680
<< metal5 >>
rect -239 7304 81 7470
rect 2221 7379 2541 7470
rect -1943 7280 1785 7304
rect -1943 2680 -1919 7280
rect 1761 2680 1785 7280
rect -1943 2656 1785 2680
rect -239 2324 81 2656
rect 2221 2581 2263 7379
rect 2499 2581 2541 7379
rect 2221 2399 2541 2581
rect -1943 2300 1785 2324
rect -1943 -2300 -1919 2300
rect 1761 -2300 1785 2300
rect -1943 -2324 1785 -2300
rect -239 -2656 81 -2324
rect 2221 -2399 2263 2399
rect 2499 -2399 2541 2399
rect 2221 -2581 2541 -2399
rect -1943 -2680 1785 -2656
rect -1943 -7280 -1919 -2680
rect 1761 -7280 1785 -2680
rect -1943 -7304 1785 -7280
rect -239 -7470 81 -7304
rect 2221 -7379 2263 -2581
rect 2499 -7379 2541 -2581
rect 2221 -7470 2541 -7379
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2519 2540 2361 7420
string parameters w 23.4 l 23.4 val 1.112k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
