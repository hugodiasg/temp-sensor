magic
tech sky130A
magscale 1 2
timestamp 1646428335
<< metal4 >>
rect -2472 7238 2472 7279
rect -2472 2534 2216 7238
rect 2452 2534 2472 7238
rect -2472 2493 2472 2534
rect -2472 2352 2472 2393
rect -2472 -2352 2216 2352
rect 2452 -2352 2472 2352
rect -2472 -2393 2472 -2352
rect -2472 -2534 2472 -2493
rect -2472 -7238 2216 -2534
rect 2452 -7238 2472 -2534
rect -2472 -7279 2472 -7238
<< via4 >>
rect 2216 2534 2452 7238
rect 2216 -2352 2452 2352
rect 2216 -7238 2452 -2534
<< mimcap2 >>
rect -2372 7139 2214 7179
rect -2372 2633 -1881 7139
rect 1723 2633 2214 7139
rect -2372 2593 2214 2633
rect -2372 2253 2214 2293
rect -2372 -2253 -1881 2253
rect 1723 -2253 2214 2253
rect -2372 -2293 2214 -2253
rect -2372 -2633 2214 -2593
rect -2372 -7139 -1881 -2633
rect 1723 -7139 2214 -2633
rect -2372 -7179 2214 -7139
<< mimcap2contact >>
rect -1881 2633 1723 7139
rect -1881 -2253 1723 2253
rect -1881 -7139 1723 -2633
<< metal5 >>
rect -239 7163 81 7329
rect 2174 7238 2494 7329
rect -1905 7139 1747 7163
rect -1905 2633 -1881 7139
rect 1723 2633 1747 7139
rect -1905 2609 1747 2633
rect -239 2277 81 2609
rect 2174 2534 2216 7238
rect 2452 2534 2494 7238
rect 2174 2352 2494 2534
rect -1905 2253 1747 2277
rect -1905 -2253 -1881 2253
rect 1723 -2253 1747 2253
rect -1905 -2277 1747 -2253
rect -239 -2609 81 -2277
rect 2174 -2352 2216 2352
rect 2452 -2352 2494 2352
rect 2174 -2534 2494 -2352
rect -1905 -2633 1747 -2609
rect -1905 -7139 -1881 -2633
rect 1723 -7139 1747 -2633
rect -1905 -7163 1747 -7139
rect -239 -7329 81 -7163
rect 2174 -7238 2216 -2534
rect 2452 -7238 2494 -2534
rect 2174 -7329 2494 -7238
<< properties >>
string FIXED_BBOX -2472 2493 2314 7279
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 22.93 l 22.93 val 1.068k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
