magic
tech sky130A
magscale 1 2
timestamp 1646019513
<< metal4 >>
rect -2662 10441 2662 10482
rect -2662 5357 2406 10441
rect 2642 5357 2662 10441
rect -2662 5316 2662 5357
rect -2662 5175 2662 5216
rect -2662 91 2406 5175
rect 2642 91 2662 5175
rect -2662 50 2662 91
rect -2662 -91 2662 -50
rect -2662 -5175 2406 -91
rect 2642 -5175 2662 -91
rect -2662 -5216 2662 -5175
rect -2662 -5357 2662 -5316
rect -2662 -10441 2406 -5357
rect 2642 -10441 2662 -5357
rect -2662 -10482 2662 -10441
<< via4 >>
rect 2406 5357 2642 10441
rect 2406 91 2642 5175
rect 2406 -5175 2642 -91
rect 2406 -10441 2642 -5357
<< mimcap2 >>
rect -2562 10342 2404 10382
rect -2562 5456 -2033 10342
rect 1875 5456 2404 10342
rect -2562 5416 2404 5456
rect -2562 5076 2404 5116
rect -2562 190 -2033 5076
rect 1875 190 2404 5076
rect -2562 150 2404 190
rect -2562 -190 2404 -150
rect -2562 -5076 -2033 -190
rect 1875 -5076 2404 -190
rect -2562 -5116 2404 -5076
rect -2562 -5456 2404 -5416
rect -2562 -10342 -2033 -5456
rect 1875 -10342 2404 -5456
rect -2562 -10382 2404 -10342
<< mimcap2contact >>
rect -2033 5456 1875 10342
rect -2033 190 1875 5076
rect -2033 -5076 1875 -190
rect -2033 -10342 1875 -5456
<< metal5 >>
rect -239 10366 81 10532
rect 2364 10441 2684 10532
rect -2057 10342 1899 10366
rect -2057 5456 -2033 10342
rect 1875 5456 1899 10342
rect -2057 5432 1899 5456
rect -239 5100 81 5432
rect 2364 5357 2406 10441
rect 2642 5357 2684 10441
rect 2364 5175 2684 5357
rect -2057 5076 1899 5100
rect -2057 190 -2033 5076
rect 1875 190 1899 5076
rect -2057 166 1899 190
rect -239 -166 81 166
rect 2364 91 2406 5175
rect 2642 91 2684 5175
rect 2364 -91 2684 91
rect -2057 -190 1899 -166
rect -2057 -5076 -2033 -190
rect 1875 -5076 1899 -190
rect -2057 -5100 1899 -5076
rect -239 -5432 81 -5100
rect 2364 -5175 2406 -91
rect 2642 -5175 2684 -91
rect 2364 -5357 2684 -5175
rect -2057 -5456 1899 -5432
rect -2057 -10342 -2033 -5456
rect 1875 -10342 1899 -5456
rect -2057 -10366 1899 -10342
rect -239 -10532 81 -10366
rect 2364 -10441 2406 -5357
rect 2642 -10441 2684 -5357
rect 2364 -10532 2684 -10441
<< properties >>
string FIXED_BBOX -2662 5316 2504 10482
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.83 l 24.83 val 1.251k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
