magic
tech sky130A
magscale 1 2
timestamp 1692041398
<< nwell >>
rect 14120 4300 14712 4938
rect 19600 4300 20192 4938
rect 14120 3400 14712 4038
rect 19600 3400 20192 4038
<< pwell >>
rect 15300 2560 15892 3180
rect 21440 2560 22032 3180
rect 14360 1680 14952 2300
rect 21440 1680 22032 2300
<< nmos >>
rect 15496 2770 15696 2970
rect 21636 2770 21836 2970
rect 14556 1890 14756 2090
rect 21636 1890 21836 2090
<< pmos >>
rect 14316 4519 14516 4719
rect 19796 4519 19996 4719
rect 14316 3619 14516 3819
rect 19796 3619 19996 3819
<< ndiff >>
rect 15438 2958 15496 2970
rect 15438 2782 15450 2958
rect 15484 2782 15496 2958
rect 15438 2770 15496 2782
rect 15696 2958 15754 2970
rect 15696 2782 15708 2958
rect 15742 2782 15754 2958
rect 15696 2770 15754 2782
rect 21578 2958 21636 2970
rect 21578 2782 21590 2958
rect 21624 2782 21636 2958
rect 21578 2770 21636 2782
rect 21836 2958 21894 2970
rect 21836 2782 21848 2958
rect 21882 2782 21894 2958
rect 21836 2770 21894 2782
rect 14498 2078 14556 2090
rect 14498 1902 14510 2078
rect 14544 1902 14556 2078
rect 14498 1890 14556 1902
rect 14756 2078 14814 2090
rect 14756 1902 14768 2078
rect 14802 1902 14814 2078
rect 14756 1890 14814 1902
rect 21578 2078 21636 2090
rect 21578 1902 21590 2078
rect 21624 1902 21636 2078
rect 21578 1890 21636 1902
rect 21836 2078 21894 2090
rect 21836 1902 21848 2078
rect 21882 1902 21894 2078
rect 21836 1890 21894 1902
<< pdiff >>
rect 14258 4707 14316 4719
rect 14258 4531 14270 4707
rect 14304 4531 14316 4707
rect 14258 4519 14316 4531
rect 14516 4707 14574 4719
rect 14516 4531 14528 4707
rect 14562 4531 14574 4707
rect 14516 4519 14574 4531
rect 19738 4707 19796 4719
rect 19738 4531 19750 4707
rect 19784 4531 19796 4707
rect 19738 4519 19796 4531
rect 19996 4707 20054 4719
rect 19996 4531 20008 4707
rect 20042 4531 20054 4707
rect 19996 4519 20054 4531
rect 14258 3807 14316 3819
rect 14258 3631 14270 3807
rect 14304 3631 14316 3807
rect 14258 3619 14316 3631
rect 14516 3807 14574 3819
rect 14516 3631 14528 3807
rect 14562 3631 14574 3807
rect 14516 3619 14574 3631
rect 19738 3807 19796 3819
rect 19738 3631 19750 3807
rect 19784 3631 19796 3807
rect 19738 3619 19796 3631
rect 19996 3807 20054 3819
rect 19996 3631 20008 3807
rect 20042 3631 20054 3807
rect 19996 3619 20054 3631
<< ndiffc >>
rect 15450 2782 15484 2958
rect 15708 2782 15742 2958
rect 21590 2782 21624 2958
rect 21848 2782 21882 2958
rect 14510 1902 14544 2078
rect 14768 1902 14802 2078
rect 21590 1902 21624 2078
rect 21848 1902 21882 2078
<< pdiffc >>
rect 14270 4531 14304 4707
rect 14528 4531 14562 4707
rect 19750 4531 19784 4707
rect 20008 4531 20042 4707
rect 14270 3631 14304 3807
rect 14528 3631 14562 3807
rect 19750 3631 19784 3807
rect 20008 3631 20042 3807
<< psubdiff >>
rect 15336 3110 15432 3144
rect 15760 3110 15856 3144
rect 15336 3048 15370 3110
rect 15822 3048 15856 3110
rect 21476 3110 21572 3144
rect 21900 3110 21996 3144
rect 15336 2630 15370 2692
rect 21476 3048 21510 3110
rect 15822 2630 15856 2692
rect 21962 3048 21996 3110
rect 15336 2596 15432 2630
rect 15760 2596 15856 2630
rect 21476 2630 21510 2692
rect 21962 2630 21996 2692
rect 21476 2596 21572 2630
rect 21900 2596 21996 2630
rect 14396 2230 14492 2264
rect 14820 2230 14916 2264
rect 14396 2168 14430 2230
rect 14882 2168 14916 2230
rect 14396 1750 14430 1812
rect 21476 2230 21572 2264
rect 21900 2230 21996 2264
rect 21476 2168 21510 2230
rect 14882 1750 14916 1812
rect 21962 2168 21996 2230
rect 14396 1716 14492 1750
rect 14820 1716 14916 1750
rect 21476 1750 21510 1812
rect 21962 1750 21996 1812
rect 21476 1716 21572 1750
rect 21900 1716 21996 1750
<< nsubdiff >>
rect 14156 4868 14252 4902
rect 14580 4868 14676 4902
rect 14156 4806 14190 4868
rect 14642 4806 14676 4868
rect 14156 4370 14190 4432
rect 14642 4370 14676 4432
rect 14156 4336 14252 4370
rect 14580 4336 14676 4370
rect 19636 4868 19732 4902
rect 20060 4868 20156 4902
rect 19636 4806 19670 4868
rect 20122 4806 20156 4868
rect 19636 4370 19670 4432
rect 20122 4370 20156 4432
rect 19636 4336 19732 4370
rect 20060 4336 20156 4370
rect 14156 3968 14252 4002
rect 14580 3968 14676 4002
rect 14156 3906 14190 3968
rect 14642 3906 14676 3968
rect 14156 3470 14190 3532
rect 14642 3470 14676 3532
rect 14156 3436 14252 3470
rect 14580 3436 14676 3470
rect 19636 3968 19732 4002
rect 20060 3968 20156 4002
rect 19636 3906 19670 3968
rect 20122 3906 20156 3968
rect 19636 3470 19670 3532
rect 20122 3470 20156 3532
rect 19636 3436 19732 3470
rect 20060 3436 20156 3470
<< psubdiffcont >>
rect 15432 3110 15760 3144
rect 15336 2692 15370 3048
rect 21572 3110 21900 3144
rect 15822 2692 15856 3048
rect 21476 2692 21510 3048
rect 15432 2596 15760 2630
rect 21962 2692 21996 3048
rect 21572 2596 21900 2630
rect 14492 2230 14820 2264
rect 14396 1812 14430 2168
rect 14882 1812 14916 2168
rect 21572 2230 21900 2264
rect 21476 1812 21510 2168
rect 14492 1716 14820 1750
rect 21962 1812 21996 2168
rect 21572 1716 21900 1750
<< nsubdiffcont >>
rect 14252 4868 14580 4902
rect 14156 4432 14190 4806
rect 14642 4432 14676 4806
rect 14252 4336 14580 4370
rect 19732 4868 20060 4902
rect 19636 4432 19670 4806
rect 20122 4432 20156 4806
rect 19732 4336 20060 4370
rect 14252 3968 14580 4002
rect 14156 3532 14190 3906
rect 14642 3532 14676 3906
rect 14252 3436 14580 3470
rect 19732 3968 20060 4002
rect 19636 3532 19670 3906
rect 20122 3532 20156 3906
rect 19732 3436 20060 3470
<< poly >>
rect 14316 4800 14516 4816
rect 14316 4766 14332 4800
rect 14500 4766 14516 4800
rect 14316 4719 14516 4766
rect 14316 4472 14516 4519
rect 14316 4438 14332 4472
rect 14500 4438 14516 4472
rect 14316 4422 14516 4438
rect 19796 4800 19996 4816
rect 19796 4766 19812 4800
rect 19980 4766 19996 4800
rect 19796 4719 19996 4766
rect 19796 4472 19996 4519
rect 19796 4438 19812 4472
rect 19980 4438 19996 4472
rect 19796 4422 19996 4438
rect 14316 3900 14516 3916
rect 14316 3866 14332 3900
rect 14500 3866 14516 3900
rect 14316 3819 14516 3866
rect 14316 3572 14516 3619
rect 14316 3538 14332 3572
rect 14500 3538 14516 3572
rect 14316 3522 14516 3538
rect 19796 3900 19996 3916
rect 19796 3866 19812 3900
rect 19980 3866 19996 3900
rect 19796 3819 19996 3866
rect 19796 3572 19996 3619
rect 19796 3538 19812 3572
rect 19980 3538 19996 3572
rect 19796 3522 19996 3538
rect 15496 3042 15696 3058
rect 15496 3008 15512 3042
rect 15680 3008 15696 3042
rect 15496 2970 15696 3008
rect 15496 2732 15696 2770
rect 15496 2698 15512 2732
rect 15680 2698 15696 2732
rect 15496 2682 15696 2698
rect 16420 3000 16730 3050
rect 17520 2990 17730 3040
rect 18570 2990 18740 3040
rect 19600 2990 19810 3050
rect 20630 3000 20900 3050
rect 16930 2690 17330 2750
rect 17990 2690 18310 2740
rect 18990 2690 19390 2740
rect 20030 2690 20430 2740
rect 21636 3042 21836 3058
rect 21636 3008 21652 3042
rect 21820 3008 21836 3042
rect 21636 2970 21836 3008
rect 21636 2732 21836 2770
rect 21636 2698 21652 2732
rect 21820 2698 21836 2732
rect 21636 2682 21836 2698
rect 14556 2162 14756 2178
rect 14556 2128 14572 2162
rect 14740 2128 14756 2162
rect 14556 2090 14756 2128
rect 14556 1852 14756 1890
rect 14556 1818 14572 1852
rect 14740 1818 14756 1852
rect 14556 1802 14756 1818
rect 16120 1800 21210 1850
rect 21636 2162 21836 2178
rect 21636 2128 21652 2162
rect 21820 2128 21836 2162
rect 21636 2090 21836 2128
rect 21636 1852 21836 1890
rect 21636 1818 21652 1852
rect 21820 1818 21836 1852
rect 21636 1802 21836 1818
<< polycont >>
rect 14332 4766 14500 4800
rect 14332 4438 14500 4472
rect 19812 4766 19980 4800
rect 19812 4438 19980 4472
rect 14332 3866 14500 3900
rect 14332 3538 14500 3572
rect 19812 3866 19980 3900
rect 19812 3538 19980 3572
rect 15512 3008 15680 3042
rect 15512 2698 15680 2732
rect 21652 3008 21820 3042
rect 21652 2698 21820 2732
rect 14572 2128 14740 2162
rect 14572 1818 14740 1852
rect 21652 2128 21820 2162
rect 21652 1818 21820 1852
<< locali >>
rect 14156 4868 14252 4902
rect 14580 4868 14676 4902
rect 14156 4806 14190 4868
rect 14642 4806 14676 4868
rect 14316 4766 14332 4800
rect 14500 4766 14516 4800
rect 14270 4707 14304 4723
rect 14270 4515 14304 4531
rect 14528 4707 14562 4723
rect 14528 4515 14562 4531
rect 14316 4438 14332 4472
rect 14500 4438 14516 4472
rect 14156 4370 14190 4432
rect 14642 4370 14676 4432
rect 14156 4336 14252 4370
rect 14580 4336 14676 4370
rect 19636 4868 19732 4902
rect 20060 4868 20156 4902
rect 19636 4806 19670 4868
rect 20122 4806 20156 4868
rect 19796 4766 19812 4800
rect 19980 4766 19996 4800
rect 19750 4707 19784 4723
rect 19750 4515 19784 4531
rect 20008 4707 20042 4723
rect 20008 4515 20042 4531
rect 19796 4438 19812 4472
rect 19980 4438 19996 4472
rect 19636 4370 19670 4432
rect 20122 4370 20156 4432
rect 19636 4336 19732 4370
rect 20060 4336 20156 4370
rect 14156 3968 14252 4002
rect 14580 3968 14676 4002
rect 14156 3906 14190 3968
rect 14642 3906 14676 3968
rect 14316 3866 14332 3900
rect 14500 3866 14516 3900
rect 14270 3807 14304 3823
rect 14270 3615 14304 3631
rect 14528 3807 14562 3823
rect 14528 3615 14562 3631
rect 14316 3538 14332 3572
rect 14500 3538 14516 3572
rect 14156 3470 14190 3532
rect 14642 3470 14676 3532
rect 14156 3436 14252 3470
rect 14580 3436 14676 3470
rect 19636 3968 19732 4002
rect 20060 3968 20156 4002
rect 19636 3906 19670 3968
rect 20122 3906 20156 3968
rect 19796 3866 19812 3900
rect 19980 3866 19996 3900
rect 19750 3807 19784 3823
rect 19750 3615 19784 3631
rect 20008 3807 20042 3823
rect 20008 3615 20042 3631
rect 19796 3538 19812 3572
rect 19980 3538 19996 3572
rect 19636 3470 19670 3532
rect 20122 3470 20156 3532
rect 19636 3436 19732 3470
rect 20060 3436 20156 3470
rect 15336 3110 15432 3144
rect 15760 3110 15856 3144
rect 15336 3048 15370 3110
rect 15822 3048 15856 3110
rect 15496 3008 15512 3042
rect 15680 3008 15696 3042
rect 15450 2958 15484 2974
rect 15450 2766 15484 2782
rect 15708 2958 15742 2974
rect 15708 2766 15742 2782
rect 15496 2698 15512 2732
rect 15680 2698 15696 2732
rect 15336 2630 15370 2692
rect 15822 2630 15856 2692
rect 15336 2596 15432 2630
rect 15760 2596 15856 2630
rect 21476 3110 21572 3144
rect 21900 3110 21996 3144
rect 21476 3048 21510 3110
rect 21962 3048 21996 3110
rect 21636 3008 21652 3042
rect 21820 3008 21836 3042
rect 21590 2958 21624 2974
rect 21590 2766 21624 2782
rect 21848 2958 21882 2974
rect 21848 2766 21882 2782
rect 21636 2698 21652 2732
rect 21820 2698 21836 2732
rect 21476 2630 21510 2692
rect 21962 2630 21996 2692
rect 21476 2596 21572 2630
rect 21900 2596 21996 2630
rect 14396 2230 14492 2264
rect 14820 2230 14916 2264
rect 14396 2168 14430 2230
rect 14882 2168 14916 2230
rect 14556 2128 14572 2162
rect 14740 2128 14756 2162
rect 14510 2078 14544 2094
rect 14510 1886 14544 1902
rect 14768 2078 14802 2094
rect 14768 1886 14802 1902
rect 14556 1818 14572 1852
rect 14740 1818 14756 1852
rect 14396 1750 14430 1812
rect 14882 1750 14916 1812
rect 14396 1716 14492 1750
rect 14820 1716 14916 1750
rect 21476 2230 21572 2264
rect 21900 2230 21996 2264
rect 21476 2168 21510 2230
rect 21962 2168 21996 2230
rect 21636 2128 21652 2162
rect 21820 2128 21836 2162
rect 21590 2078 21624 2094
rect 21590 1886 21624 1902
rect 21848 2078 21882 2094
rect 21848 1886 21882 1902
rect 21636 1818 21652 1852
rect 21820 1818 21836 1852
rect 21476 1750 21510 1812
rect 21962 1750 21996 1812
rect 21476 1716 21572 1750
rect 21900 1716 21996 1750
<< metal1 >>
rect 15160 4780 19150 4830
rect 15110 4700 16935 4730
rect 15110 4240 15150 4700
rect 16610 4590 16690 4600
rect 16610 4580 16620 4590
rect 15380 4550 16620 4580
rect 16610 4520 16620 4550
rect 16680 4520 16690 4590
rect 16610 4510 16690 4520
rect 16980 4240 17020 4720
rect 17280 4410 17330 4780
rect 18110 4700 19380 4730
rect 17620 4590 17700 4600
rect 17620 4520 17630 4590
rect 17690 4580 17700 4590
rect 17690 4550 19110 4580
rect 17690 4520 17700 4550
rect 17620 4510 17700 4520
rect 17280 4400 17360 4410
rect 17280 4340 17290 4400
rect 17350 4340 17360 4400
rect 17280 4330 17360 4340
rect 17280 4300 17330 4330
rect 19260 4240 19380 4700
rect 13875 4110 19380 4240
rect 15110 3830 15150 4110
rect 15110 3800 16935 3830
rect 16610 3710 16710 3720
rect 16610 3680 16620 3710
rect 15380 3650 16620 3680
rect 16610 3620 16620 3650
rect 16700 3620 16710 3710
rect 16610 3610 16710 3620
rect 16980 3610 17020 4110
rect 19260 3830 19380 4110
rect 17280 3570 17310 3820
rect 18120 3800 19380 3830
rect 19260 3760 19380 3800
rect 17580 3710 17680 3720
rect 17580 3620 17590 3710
rect 17670 3680 17680 3710
rect 17670 3650 18940 3680
rect 17670 3620 17680 3650
rect 17580 3610 17680 3620
rect 15170 3520 19140 3570
rect 17280 3385 17310 3520
rect 17280 3355 17635 3385
rect 13880 3230 13990 3270
rect 13880 3190 15660 3230
rect 17605 3210 17635 3355
rect 13880 3160 13990 3190
rect 15620 2730 15660 3190
rect 16060 3170 21270 3210
rect 16060 2880 16100 3170
rect 16320 3080 16880 3120
rect 16170 2730 16180 2770
rect 15620 2700 16180 2730
rect 16270 2700 16280 2770
rect 15620 2690 16280 2700
rect 16320 2660 16360 3080
rect 16680 3040 16790 3050
rect 16680 2960 16690 3040
rect 16780 2960 16790 3040
rect 16680 2950 16790 2960
rect 15650 2620 16360 2660
rect 13880 2340 13990 2380
rect 13880 2300 15160 2340
rect 13880 2270 13990 2300
rect 15120 2160 15160 2300
rect 15120 2120 15620 2160
rect 15120 1920 15160 2120
rect 15380 1680 15420 2040
rect 15650 1900 15690 2620
rect 16575 2575 16625 2905
rect 16840 2660 16880 3080
rect 17100 2890 17140 3170
rect 17360 3080 17920 3120
rect 16920 2770 17030 2780
rect 16920 2700 16930 2770
rect 17020 2700 17030 2770
rect 16920 2690 17030 2700
rect 17180 2770 17300 2780
rect 17180 2700 17190 2770
rect 17290 2700 17300 2770
rect 17180 2690 17300 2700
rect 17360 2660 17400 3080
rect 17450 3040 17560 3050
rect 17450 2960 17460 3040
rect 17550 2960 17560 3040
rect 17450 2950 17560 2960
rect 17710 3040 17820 3050
rect 17710 2960 17720 3040
rect 17810 2960 17820 3040
rect 17710 2950 17820 2960
rect 16840 2620 17400 2660
rect 17605 2590 17655 2905
rect 17880 2660 17920 3080
rect 18130 2890 18170 3170
rect 18390 3080 18940 3120
rect 17950 2770 18070 2780
rect 17950 2700 17960 2770
rect 18060 2700 18070 2770
rect 17950 2690 18070 2700
rect 18220 2770 18340 2780
rect 18220 2700 18230 2770
rect 18330 2700 18340 2770
rect 18220 2690 18340 2700
rect 18390 2660 18430 3080
rect 18480 3040 18590 3050
rect 18480 2960 18490 3040
rect 18580 2960 18590 3040
rect 18480 2950 18590 2960
rect 18740 3040 18850 3050
rect 18740 2960 18750 3040
rect 18840 2960 18850 3040
rect 18740 2950 18850 2960
rect 17880 2620 18430 2660
rect 17570 2575 17655 2590
rect 18645 2575 18695 2945
rect 18900 2660 18940 3080
rect 19160 2890 19200 3170
rect 19420 3080 19980 3120
rect 18980 2770 19100 2780
rect 18980 2700 18990 2770
rect 19090 2700 19100 2770
rect 18980 2690 19100 2700
rect 19250 2770 19370 2780
rect 19250 2700 19260 2770
rect 19360 2700 19370 2770
rect 19250 2690 19370 2700
rect 19420 2660 19460 3080
rect 19520 3030 19630 3040
rect 19520 2950 19530 3030
rect 19620 2950 19630 3030
rect 19520 2940 19630 2950
rect 19770 3030 19880 3040
rect 19770 2950 19780 3030
rect 19870 2950 19880 3030
rect 19770 2940 19880 2950
rect 18900 2620 19460 2660
rect 19675 2575 19725 2905
rect 19940 2660 19980 3080
rect 20200 2890 20240 3170
rect 20450 3080 21010 3120
rect 20020 2770 20140 2780
rect 20020 2700 20030 2770
rect 20130 2700 20140 2770
rect 20020 2690 20140 2700
rect 20270 2770 20390 2780
rect 20270 2700 20280 2770
rect 20380 2700 20390 2770
rect 20270 2690 20390 2700
rect 20450 2660 20490 3080
rect 20540 3030 20650 3040
rect 20540 2950 20550 3030
rect 20640 2950 20650 3030
rect 20540 2940 20650 2950
rect 19940 2620 20490 2660
rect 20705 2575 20755 2905
rect 20970 2880 21010 3080
rect 21230 2900 21270 3170
rect 21050 2760 21170 2770
rect 16570 2560 20755 2575
rect 16570 2525 17270 2560
rect 17260 2480 17270 2525
rect 17370 2525 20755 2560
rect 20840 2530 20880 2730
rect 21050 2690 21060 2760
rect 21160 2690 21170 2760
rect 21050 2680 21170 2690
rect 17370 2480 17380 2525
rect 17570 2510 17650 2525
rect 20840 2490 21420 2530
rect 17100 2470 17200 2480
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 21380 2340 21420 2490
rect 16840 2300 22120 2340
rect 16060 2210 16620 2250
rect 16060 1680 16100 2210
rect 16130 1856 16180 1860
rect 16130 1850 16258 1856
rect 16320 1850 16360 2080
rect 16130 1820 16360 1850
rect 16150 1810 16360 1820
rect 15380 1640 16100 1680
rect 15710 1430 16100 1640
rect 16168 1520 16258 1810
rect 16320 1680 16360 1810
rect 16580 1780 16620 2210
rect 16840 1950 16880 2300
rect 17100 2210 17660 2250
rect 17100 1780 17140 2210
rect 16580 1740 17140 1780
rect 17100 1708 17200 1710
rect 17100 1680 17113 1708
rect 16320 1640 17113 1680
rect 17100 1633 17113 1640
rect 17188 1680 17200 1708
rect 17360 1680 17400 1960
rect 17620 1780 17660 2210
rect 17870 1970 17910 2300
rect 18130 2210 18690 2250
rect 18130 1780 18170 2210
rect 17620 1740 18170 1780
rect 18390 1680 18430 1970
rect 18650 1770 18690 2210
rect 18900 1950 18940 2300
rect 19160 2210 19720 2250
rect 19160 1770 19200 2210
rect 18650 1730 19200 1770
rect 19420 1680 19460 1960
rect 19680 1780 19720 2210
rect 19940 1960 19980 2300
rect 20190 2210 20750 2250
rect 20190 1780 20230 2210
rect 19680 1740 20230 1780
rect 20450 1680 20490 1960
rect 20710 1780 20750 2210
rect 20970 1950 21010 2300
rect 21230 1780 21270 2000
rect 20710 1740 21270 1780
rect 17188 1640 20490 1680
rect 17188 1633 17200 1640
rect 17100 1620 17200 1633
rect 17844 1540 18090 1542
rect 17840 1532 18090 1540
rect 17134 1520 17380 1522
rect 16168 1512 17380 1520
rect 16168 1430 17146 1512
rect 17134 1252 17146 1430
rect 17364 1252 17380 1512
rect 17840 1450 17856 1532
rect 17844 1272 17856 1450
rect 18074 1503 18090 1532
rect 18074 1500 18190 1503
rect 22010 1500 22120 2300
rect 18074 1393 22120 1500
rect 18074 1272 18090 1393
rect 18190 1390 22120 1393
rect 17844 1260 18090 1272
rect 17134 1238 17380 1252
<< via1 >>
rect 16620 4520 16680 4590
rect 17630 4520 17690 4590
rect 17290 4340 17350 4400
rect 16620 3620 16700 3710
rect 17590 3620 17670 3710
rect 16180 2700 16270 2770
rect 16690 2960 16780 3040
rect 16930 2700 17020 2770
rect 17190 2700 17290 2770
rect 17460 2960 17550 3040
rect 17720 2960 17810 3040
rect 17960 2700 18060 2770
rect 18230 2700 18330 2770
rect 18490 2960 18580 3040
rect 18750 2960 18840 3040
rect 18990 2700 19090 2770
rect 19260 2700 19360 2770
rect 19530 2950 19620 3030
rect 19780 2950 19870 3030
rect 20030 2700 20130 2770
rect 20280 2700 20380 2770
rect 20550 2950 20640 3030
rect 17270 2480 17370 2560
rect 21060 2690 21160 2760
rect 17110 2390 17190 2470
rect 17113 1633 17188 1708
rect 17146 1252 17364 1512
rect 17856 1272 18074 1532
<< metal2 >>
rect 16610 4590 16690 4600
rect 16610 4520 16620 4590
rect 16680 4520 16690 4590
rect 16610 4510 16690 4520
rect 17620 4590 17700 4600
rect 17620 4520 17630 4590
rect 17690 4520 17700 4590
rect 17620 4510 17700 4520
rect 17280 4400 17360 4410
rect 17280 4340 17290 4400
rect 17350 4340 17360 4400
rect 16610 3710 16710 3720
rect 16610 3620 16620 3710
rect 16700 3620 16710 3710
rect 16610 3460 16710 3620
rect 16610 3360 16780 3460
rect 16680 3050 16780 3360
rect 17280 3330 17360 4340
rect 17405 3710 17680 3720
rect 17405 3620 17590 3710
rect 17670 3620 17680 3710
rect 17405 3610 17680 3620
rect 17270 3320 17370 3330
rect 17270 3230 17370 3240
rect 17405 3050 17515 3610
rect 16680 3040 17560 3050
rect 16680 2960 16690 3040
rect 16780 2960 17460 3040
rect 17550 2960 17560 3040
rect 16680 2950 17560 2960
rect 17710 3040 18590 3050
rect 17710 2960 17720 3040
rect 17810 2960 18490 3040
rect 18580 2960 18590 3040
rect 17710 2950 18590 2960
rect 18740 3040 19630 3050
rect 18740 2960 18750 3040
rect 18840 3030 19630 3040
rect 18840 2960 19530 3030
rect 18740 2950 19530 2960
rect 19620 2950 19630 3030
rect 18740 2940 19630 2950
rect 19770 3030 20650 3040
rect 19770 2950 19780 3030
rect 19870 2950 20550 3030
rect 20640 2950 20650 3030
rect 19770 2940 19880 2950
rect 20540 2940 20650 2950
rect 16180 2770 16270 2780
rect 16170 2700 16180 2760
rect 16920 2770 17030 2780
rect 16270 2740 16280 2760
rect 16920 2740 16930 2770
rect 16270 2700 16930 2740
rect 17020 2740 17030 2770
rect 17180 2770 17300 2780
rect 17020 2700 17040 2740
rect 16170 2690 17040 2700
rect 17180 2700 17190 2770
rect 17290 2700 17300 2770
rect 17180 2690 17300 2700
rect 17950 2770 18070 2780
rect 17950 2700 17960 2770
rect 18060 2700 18070 2770
rect 17950 2690 18070 2700
rect 18220 2770 19100 2780
rect 18220 2700 18230 2770
rect 18330 2700 18990 2770
rect 19090 2700 19100 2770
rect 18220 2690 19100 2700
rect 19250 2770 20140 2780
rect 19250 2700 19260 2770
rect 19360 2700 20030 2770
rect 20130 2700 20140 2770
rect 19250 2690 20140 2700
rect 20270 2770 21150 2780
rect 20270 2700 20280 2770
rect 20380 2760 21170 2770
rect 20380 2700 21060 2760
rect 20270 2690 21060 2700
rect 21160 2690 21170 2760
rect 21050 2680 21170 2690
rect 17260 2560 17380 2570
rect 17260 2480 17270 2560
rect 17370 2480 17380 2560
rect 17100 2470 17200 2480
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 17113 1710 17188 1718
rect 17100 1708 17200 1710
rect 17100 1633 17113 1708
rect 17188 1633 17200 1708
rect 17100 1620 17200 1633
rect 17844 1532 18090 1542
rect 17134 1512 17380 1522
rect 17134 1252 17146 1512
rect 17364 1252 17380 1512
rect 17844 1272 17856 1532
rect 18074 1272 18090 1532
rect 17844 1260 18090 1272
rect 17134 1238 17380 1252
<< via2 >>
rect 16620 4520 16680 4590
rect 17630 4520 17690 4590
rect 17270 3240 17370 3320
rect 17190 2700 17290 2770
rect 17960 2700 18060 2770
rect 17270 2480 17370 2560
rect 17110 2390 17190 2470
rect 17113 1633 17188 1708
rect 17146 1252 17364 1512
rect 17856 1272 18074 1532
<< metal3 >>
rect 16610 4590 17700 4600
rect 16610 4520 16620 4590
rect 16680 4520 17630 4590
rect 17690 4520 17700 4590
rect 16610 4510 17700 4520
rect 17110 3610 17190 4510
rect 17113 3390 17188 3610
rect 17100 3310 17110 3390
rect 17190 3310 17200 3390
rect 17260 3320 17380 3330
rect 17260 3240 17270 3320
rect 17370 3240 17380 3320
rect 17260 3230 17380 3240
rect 17180 2770 18070 2780
rect 17180 2700 17190 2770
rect 17290 2700 17960 2770
rect 18060 2700 18070 2770
rect 17180 2680 18070 2700
rect 17260 2560 17380 2570
rect 17113 2480 17188 2500
rect 17260 2480 17270 2560
rect 17370 2480 17380 2560
rect 17100 2470 17200 2480
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 17113 1713 17188 2380
rect 17103 1710 17198 1713
rect 17100 1708 17200 1710
rect 17100 1633 17113 1708
rect 17188 1633 17200 1708
rect 17100 1620 17200 1633
rect 17844 1532 18090 1542
rect 17134 1512 17380 1522
rect 17134 1252 17146 1512
rect 17364 1252 17380 1512
rect 17844 1272 17856 1532
rect 18074 1272 18090 1532
rect 17844 1260 18090 1272
rect 17134 1238 17380 1252
<< via3 >>
rect 17110 3310 17190 3390
rect 17270 3240 17370 3320
rect 17270 2480 17370 2560
rect 17110 2390 17190 2470
rect 17146 1252 17364 1512
rect 17856 1272 18074 1532
<< metal4 >>
rect 17101 3390 17199 3399
rect 17100 3310 17110 3390
rect 17190 3310 17200 3390
rect 17100 3300 17200 3310
rect 17260 3320 17380 3340
rect 17101 2520 17199 3300
rect 17260 3240 17270 3320
rect 17370 3240 17380 3320
rect 17260 2560 17380 3240
rect 17100 2470 17200 2520
rect 17260 2480 17270 2560
rect 17370 2480 17380 2560
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 17830 1532 18190 1580
rect 17134 1512 17380 1522
rect 17134 1384 17146 1512
rect 17130 1252 17146 1384
rect 17364 1252 17380 1512
rect 17130 928 17380 1252
rect 17830 1272 17856 1532
rect 18074 1530 18190 1532
rect 18160 1280 18190 1530
rect 18074 1272 18190 1280
rect 17830 1240 18190 1272
<< via4 >>
rect 17860 1280 18074 1530
rect 18074 1280 18160 1530
<< metal5 >>
rect 17830 1530 18190 1580
rect 17830 1280 17860 1530
rect 18160 1280 18190 1530
rect 17830 890 18190 1280
<< comment >>
rect 15530 4550 15940 4700
rect 17080 4540 17220 4700
rect 18220 4560 18630 4710
rect 15490 3640 15900 3790
rect 17100 3620 17240 3780
rect 18400 3630 18810 3780
rect 17940 2800 18620 2940
rect 15150 1910 15640 2070
rect 17940 1920 18620 2060
use sky130_fd_pr__cap_mim_m3_2_ZFPS3R  sky130_fd_pr__cap_mim_m3_2_ZFPS3R_0
timestamp 1692040603
transform 1 0 18733 0 1 -1023
box -2449 -2181 2471 2181
use sky130_fd_pr__nfet_01v8_CL66SD  sky130_fd_pr__nfet_01v8_CL66SD_0
timestamp 1661536226
transform 1 0 18667 0 1 2870
box -2747 -310 2747 310
use sky130_fd_pr__nfet_01v8_CL66SD  sky130_fd_pr__nfet_01v8_CL66SD_1
timestamp 1661536226
transform 1 0 18667 0 1 1990
box -2747 -310 2747 310
use sky130_fd_pr__nfet_01v8_GVTB53  sky130_fd_pr__nfet_01v8_GVTB53_0
timestamp 1661301161
transform 1 0 15405 0 1 1990
box -425 -310 425 310
use sky130_fd_pr__pfet_01v8_8C4HA7  sky130_fd_pr__pfet_01v8_8C4HA7_0
timestamp 1661301161
transform 1 0 15792 0 1 3719
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_8L4H97  sky130_fd_pr__pfet_01v8_8L4H97_1
timestamp 1661301161
transform 1 0 15792 0 1 4619
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_8LYGA7  sky130_fd_pr__pfet_01v8_8LYGA7_0
timestamp 1661301161
transform -1 0 18532 0 1 4619
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_8LYGA7  sky130_fd_pr__pfet_01v8_8LYGA7_1
timestamp 1661301161
transform -1 0 18532 0 1 3719
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_BLSBYX  sky130_fd_pr__pfet_01v8_BLSBYX_1
timestamp 1661301161
transform 1 0 17156 0 1 3719
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_BLSBYX  sky130_fd_pr__pfet_01v8_BLSBYX_2
timestamp 1661301161
transform 1 0 17156 0 1 4619
box -296 -319 296 319
<< labels >>
flabel metal1 19710 1650 19750 1660 0 FreeSans 800 0 0 0 net1
flabel metal1 15710 1490 15820 1600 0 FreeSans 1600 0 0 0 gnd
port 4 nsew
flabel comment 15220 1920 15340 2050 0 FreeSans 800 0 0 0 M10
flabel comment 15470 1920 15590 2050 0 FreeSans 800 0 0 0 M5
flabel comment 15490 3640 15900 3790 0 FreeSans 800 0 0 0 M6_1
flabel comment 18220 4560 18630 4710 0 FreeSans 800 0 0 0 M8_2
flabel comment 15530 4550 15940 4700 0 FreeSans 800 0 0 0 M8_1
flabel comment 17080 4540 17220 4700 0 FreeSans 800 0 0 0 M3
flabel comment 18400 3630 18810 3780 0 FreeSans 800 0 0 0 M6_2
flabel metal2 17320 4070 17320 4070 0 FreeSans 800 0 0 0 net2
flabel comment 17100 3620 17240 3780 0 FreeSans 800 0 0 0 M4
flabel metal1 15670 2390 15680 2410 0 FreeSans 800 0 0 0 net4
flabel comment 17940 1920 18620 2060 0 FreeSans 800 0 0 0 M9_M7
flabel comment 17940 2800 18620 2940 0 FreeSans 800 0 0 0 M1_M2
flabel metal1 17600 3360 17620 3380 0 FreeSans 800 0 0 0 net3
flabel metal1 13880 4120 13990 4230 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 13880 3160 13990 3270 0 FreeSans 1600 0 0 0 in
port 3 nsew
flabel metal1 13880 2270 13990 2380 0 FreeSans 1600 0 0 0 ib
port 1 nsew
flabel metal1 22010 2230 22120 2340 0 FreeSans 1600 0 0 0 out
port 2 nsew
<< end >>
