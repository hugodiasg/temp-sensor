magic
tech sky130A
magscale 1 2
timestamp 1646426843
<< metal4 >>
rect -2619 7679 2619 7720
rect -2619 2681 2363 7679
rect 2599 2681 2619 7679
rect -2619 2640 2619 2681
rect -2619 2499 2619 2540
rect -2619 -2499 2363 2499
rect 2599 -2499 2619 2499
rect -2619 -2540 2619 -2499
rect -2619 -2681 2619 -2640
rect -2619 -7679 2363 -2681
rect 2599 -7679 2619 -2681
rect -2619 -7720 2619 -7679
<< via4 >>
rect 2363 2681 2599 7679
rect 2363 -2499 2599 2499
rect 2363 -7679 2599 -2681
<< mimcap2 >>
rect -2519 7580 2361 7620
rect -2519 2780 -1999 7580
rect 1841 2780 2361 7580
rect -2519 2740 2361 2780
rect -2519 2400 2361 2440
rect -2519 -2400 -1999 2400
rect 1841 -2400 2361 2400
rect -2519 -2440 2361 -2400
rect -2519 -2780 2361 -2740
rect -2519 -7580 -1999 -2780
rect 1841 -7580 2361 -2780
rect -2519 -7620 2361 -7580
<< mimcap2contact >>
rect -1999 2780 1841 7580
rect -1999 -2400 1841 2400
rect -1999 -7580 1841 -2780
<< metal5 >>
rect -239 7604 81 7770
rect 2321 7679 2641 7770
rect -2023 7580 1865 7604
rect -2023 2780 -1999 7580
rect 1841 2780 1865 7580
rect -2023 2756 1865 2780
rect -239 2424 81 2756
rect 2321 2681 2363 7679
rect 2599 2681 2641 7679
rect 2321 2499 2641 2681
rect -2023 2400 1865 2424
rect -2023 -2400 -1999 2400
rect 1841 -2400 1865 2400
rect -2023 -2424 1865 -2400
rect -239 -2756 81 -2424
rect 2321 -2499 2363 2499
rect 2599 -2499 2641 2499
rect 2321 -2681 2641 -2499
rect -2023 -2780 1865 -2756
rect -2023 -7580 -1999 -2780
rect 1841 -7580 1865 -2780
rect -2023 -7604 1865 -7580
rect -239 -7770 81 -7604
rect 2321 -7679 2363 -2681
rect 2599 -7679 2641 -2681
rect 2321 -7770 2641 -7679
<< properties >>
string FIXED_BBOX -2619 2640 2461 7720
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.4 l 24.4 val 1.209k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
