magic
tech sky130A
magscale 1 2
timestamp 1645148224
<< metal4 >>
rect -2843 8351 2843 8392
rect -2843 2905 2587 8351
rect 2823 2905 2843 8351
rect -2843 2864 2843 2905
rect -2843 2723 2843 2764
rect -2843 -2723 2587 2723
rect 2823 -2723 2843 2723
rect -2843 -2764 2843 -2723
rect -2843 -2905 2843 -2864
rect -2843 -8351 2587 -2905
rect 2823 -8351 2843 -2905
rect -2843 -8392 2843 -8351
<< via4 >>
rect 2587 2905 2823 8351
rect 2587 -2723 2823 2723
rect 2587 -8351 2823 -2905
<< mimcap2 >>
rect -2743 8252 2585 8292
rect -2743 3004 -2178 8252
rect 2020 3004 2585 8252
rect -2743 2964 2585 3004
rect -2743 2624 2585 2664
rect -2743 -2624 -2178 2624
rect 2020 -2624 2585 2624
rect -2743 -2664 2585 -2624
rect -2743 -3004 2585 -2964
rect -2743 -8252 -2178 -3004
rect 2020 -8252 2585 -3004
rect -2743 -8292 2585 -8252
<< mimcap2contact >>
rect -2178 3004 2020 8252
rect -2178 -2624 2020 2624
rect -2178 -8252 2020 -3004
<< metal5 >>
rect -239 8276 81 8442
rect 2545 8351 2865 8442
rect -2202 8252 2044 8276
rect -2202 3004 -2178 8252
rect 2020 3004 2044 8252
rect -2202 2980 2044 3004
rect -239 2648 81 2980
rect 2545 2905 2587 8351
rect 2823 2905 2865 8351
rect 2545 2723 2865 2905
rect -2202 2624 2044 2648
rect -2202 -2624 -2178 2624
rect 2020 -2624 2044 2624
rect -2202 -2648 2044 -2624
rect -239 -2980 81 -2648
rect 2545 -2723 2587 2723
rect 2823 -2723 2865 2723
rect 2545 -2905 2865 -2723
rect -2202 -3004 2044 -2980
rect -2202 -8252 -2178 -3004
rect 2020 -8252 2044 -3004
rect -2202 -8276 2044 -8252
rect -239 -8442 81 -8276
rect 2545 -8351 2587 -2905
rect 2823 -8351 2865 -2905
rect 2545 -8442 2865 -8351
<< properties >>
string FIXED_BBOX -2843 2864 2685 8392
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 26.643 l 26.643 val 1.439k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
