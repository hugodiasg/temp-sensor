magic
tech sky130A
magscale 1 2
timestamp 1661709424
<< nwell >>
rect 14130 4300 14722 4938
rect 19600 4310 20192 4948
rect 14130 3400 14722 4038
rect 19600 3400 20192 4038
<< pwell >>
rect 15330 2560 15922 3180
rect 21410 2560 22002 3180
rect 14390 1680 14980 2300
rect 21420 1680 22010 2300
<< nmos >>
rect 15526 2770 15726 2970
rect 21606 2770 21806 2970
rect 14586 1890 14786 2090
rect 21616 1890 21816 2090
<< pmos >>
rect 14326 4519 14526 4719
rect 19796 4529 19996 4729
rect 14326 3619 14526 3819
rect 19796 3619 19996 3819
<< ndiff >>
rect 15468 2958 15526 2970
rect 15468 2782 15480 2958
rect 15514 2782 15526 2958
rect 15468 2770 15526 2782
rect 15726 2958 15784 2970
rect 15726 2782 15738 2958
rect 15772 2782 15784 2958
rect 15726 2770 15784 2782
rect 21548 2958 21606 2970
rect 21548 2782 21560 2958
rect 21594 2782 21606 2958
rect 21548 2770 21606 2782
rect 21806 2958 21864 2970
rect 21806 2782 21818 2958
rect 21852 2782 21864 2958
rect 21806 2770 21864 2782
rect 14528 2078 14586 2090
rect 14528 1902 14540 2078
rect 14574 1902 14586 2078
rect 14528 1890 14586 1902
rect 14786 2078 14844 2090
rect 14786 1902 14798 2078
rect 14832 1902 14844 2078
rect 14786 1890 14844 1902
rect 21558 2078 21616 2090
rect 21558 1902 21570 2078
rect 21604 1902 21616 2078
rect 21558 1890 21616 1902
rect 21816 2078 21874 2090
rect 21816 1902 21828 2078
rect 21862 1902 21874 2078
rect 21816 1890 21874 1902
<< pdiff >>
rect 14268 4707 14326 4719
rect 14268 4531 14280 4707
rect 14314 4531 14326 4707
rect 14268 4519 14326 4531
rect 14526 4707 14584 4719
rect 14526 4531 14538 4707
rect 14572 4531 14584 4707
rect 14526 4519 14584 4531
rect 19738 4717 19796 4729
rect 19738 4541 19750 4717
rect 19784 4541 19796 4717
rect 19738 4529 19796 4541
rect 19996 4717 20054 4729
rect 19996 4541 20008 4717
rect 20042 4541 20054 4717
rect 19996 4529 20054 4541
rect 14268 3807 14326 3819
rect 14268 3631 14280 3807
rect 14314 3631 14326 3807
rect 14268 3619 14326 3631
rect 14526 3807 14584 3819
rect 14526 3631 14538 3807
rect 14572 3631 14584 3807
rect 14526 3619 14584 3631
rect 19738 3807 19796 3819
rect 19738 3631 19750 3807
rect 19784 3631 19796 3807
rect 19738 3619 19796 3631
rect 19996 3807 20054 3819
rect 19996 3631 20008 3807
rect 20042 3631 20054 3807
rect 19996 3619 20054 3631
<< ndiffc >>
rect 15480 2782 15514 2958
rect 15738 2782 15772 2958
rect 21560 2782 21594 2958
rect 21818 2782 21852 2958
rect 14540 1902 14574 2078
rect 14798 1902 14832 2078
rect 21570 1902 21604 2078
rect 21828 1902 21862 2078
<< pdiffc >>
rect 14280 4531 14314 4707
rect 14538 4531 14572 4707
rect 19750 4541 19784 4717
rect 20008 4541 20042 4717
rect 14280 3631 14314 3807
rect 14538 3631 14572 3807
rect 19750 3631 19784 3807
rect 20008 3631 20042 3807
<< psubdiff >>
rect 15366 3110 15462 3144
rect 15790 3110 15886 3144
rect 15366 3048 15400 3110
rect 15852 3048 15886 3110
rect 21446 3110 21542 3144
rect 21870 3110 21966 3144
rect 15366 2630 15400 2692
rect 21446 3048 21480 3110
rect 15852 2630 15886 2692
rect 21932 3048 21966 3110
rect 15366 2596 15462 2630
rect 15790 2596 15886 2630
rect 21446 2630 21480 2692
rect 21932 2630 21966 2692
rect 21446 2596 21542 2630
rect 21870 2596 21966 2630
rect 14426 2230 14522 2264
rect 14850 2230 14946 2264
rect 14426 2168 14460 2230
rect 14912 2168 14946 2230
rect 14426 1750 14460 1812
rect 21456 2230 21552 2264
rect 21880 2230 21976 2264
rect 21456 2168 21490 2230
rect 14912 1750 14946 1812
rect 21942 2168 21976 2230
rect 14426 1716 14522 1750
rect 14850 1716 14946 1750
rect 21456 1750 21490 1812
rect 21942 1750 21976 1812
rect 21456 1716 21552 1750
rect 21880 1716 21976 1750
rect 15806 1490 15830 1630
rect 16020 1490 16044 1630
<< nsubdiff >>
rect 14166 4868 14262 4902
rect 14590 4868 14686 4902
rect 14166 4806 14200 4868
rect 14652 4806 14686 4868
rect 14166 4370 14200 4432
rect 14652 4370 14686 4432
rect 14166 4336 14262 4370
rect 14590 4336 14686 4370
rect 19636 4878 19732 4912
rect 20060 4878 20156 4912
rect 19636 4816 19670 4878
rect 20122 4816 20156 4878
rect 19636 4380 19670 4442
rect 20122 4380 20156 4442
rect 19636 4346 19732 4380
rect 20060 4346 20156 4380
rect 14166 3968 14262 4002
rect 14590 3968 14686 4002
rect 14166 3906 14200 3968
rect 14652 3906 14686 3968
rect 14166 3470 14200 3532
rect 14652 3470 14686 3532
rect 14166 3436 14262 3470
rect 14590 3436 14686 3470
rect 19636 3968 19732 4002
rect 20060 3968 20156 4002
rect 19636 3906 19670 3968
rect 20122 3906 20156 3968
rect 19636 3470 19670 3532
rect 20122 3470 20156 3532
rect 19636 3436 19732 3470
rect 20060 3436 20156 3470
<< psubdiffcont >>
rect 15462 3110 15790 3144
rect 15366 2692 15400 3048
rect 21542 3110 21870 3144
rect 15852 2692 15886 3048
rect 21446 2692 21480 3048
rect 15462 2596 15790 2630
rect 21932 2692 21966 3048
rect 21542 2596 21870 2630
rect 14522 2230 14850 2264
rect 14426 1812 14460 2168
rect 14912 1812 14946 2168
rect 21552 2230 21880 2264
rect 21456 1812 21490 2168
rect 14522 1716 14850 1750
rect 21942 1812 21976 2168
rect 21552 1716 21880 1750
rect 15830 1490 16020 1630
<< nsubdiffcont >>
rect 14262 4868 14590 4902
rect 14166 4432 14200 4806
rect 14652 4432 14686 4806
rect 14262 4336 14590 4370
rect 19732 4878 20060 4912
rect 19636 4442 19670 4816
rect 20122 4442 20156 4816
rect 19732 4346 20060 4380
rect 14262 3968 14590 4002
rect 14166 3532 14200 3906
rect 14652 3532 14686 3906
rect 14262 3436 14590 3470
rect 19732 3968 20060 4002
rect 19636 3532 19670 3906
rect 20122 3532 20156 3906
rect 19732 3436 20060 3470
<< poly >>
rect 14326 4800 14526 4816
rect 14326 4766 14342 4800
rect 14510 4766 14526 4800
rect 14326 4719 14526 4766
rect 14326 4472 14526 4519
rect 14326 4438 14342 4472
rect 14510 4438 14526 4472
rect 14326 4422 14526 4438
rect 19796 4810 19996 4826
rect 19796 4776 19812 4810
rect 19980 4776 19996 4810
rect 19796 4729 19996 4776
rect 19796 4482 19996 4529
rect 19796 4448 19812 4482
rect 19980 4448 19996 4482
rect 19796 4432 19996 4448
rect 14326 3900 14526 3916
rect 14326 3866 14342 3900
rect 14510 3866 14526 3900
rect 14326 3819 14526 3866
rect 14326 3572 14526 3619
rect 14326 3538 14342 3572
rect 14510 3538 14526 3572
rect 14326 3522 14526 3538
rect 19796 3900 19996 3916
rect 19796 3866 19812 3900
rect 19980 3866 19996 3900
rect 19796 3819 19996 3866
rect 19796 3572 19996 3619
rect 19796 3538 19812 3572
rect 19980 3538 19996 3572
rect 19796 3522 19996 3538
rect 15526 3042 15726 3058
rect 15526 3008 15542 3042
rect 15710 3008 15726 3042
rect 15526 2970 15726 3008
rect 15526 2732 15726 2770
rect 15526 2698 15542 2732
rect 15710 2698 15726 2732
rect 15526 2682 15726 2698
rect 16420 3000 16730 3050
rect 17520 2990 17730 3040
rect 18570 2990 18740 3040
rect 19600 2990 19810 3050
rect 20630 3000 20900 3050
rect 16930 2690 17330 2750
rect 17990 2690 18310 2740
rect 18990 2690 19390 2740
rect 20030 2690 20430 2740
rect 21606 3042 21806 3058
rect 21606 3008 21622 3042
rect 21790 3008 21806 3042
rect 21606 2970 21806 3008
rect 21606 2732 21806 2770
rect 21606 2698 21622 2732
rect 21790 2698 21806 2732
rect 21606 2682 21806 2698
rect 14586 2162 14786 2178
rect 14586 2128 14602 2162
rect 14770 2128 14786 2162
rect 14586 2090 14786 2128
rect 14586 1852 14786 1890
rect 14586 1818 14602 1852
rect 14770 1818 14786 1852
rect 14586 1802 14786 1818
rect 16120 1800 21210 1850
rect 21616 2162 21816 2178
rect 21616 2128 21632 2162
rect 21800 2128 21816 2162
rect 21616 2090 21816 2128
rect 21616 1852 21816 1890
rect 21616 1818 21632 1852
rect 21800 1818 21816 1852
rect 21616 1802 21816 1818
<< polycont >>
rect 14342 4766 14510 4800
rect 14342 4438 14510 4472
rect 19812 4776 19980 4810
rect 19812 4448 19980 4482
rect 14342 3866 14510 3900
rect 14342 3538 14510 3572
rect 19812 3866 19980 3900
rect 19812 3538 19980 3572
rect 15542 3008 15710 3042
rect 15542 2698 15710 2732
rect 21622 3008 21790 3042
rect 21622 2698 21790 2732
rect 14602 2128 14770 2162
rect 14602 1818 14770 1852
rect 21632 2128 21800 2162
rect 21632 1818 21800 1852
<< locali >>
rect 14166 4868 14262 4902
rect 14590 4868 14686 4902
rect 14166 4806 14200 4868
rect 14652 4806 14686 4868
rect 14326 4766 14342 4800
rect 14510 4766 14526 4800
rect 14280 4707 14314 4723
rect 14280 4515 14314 4531
rect 14538 4707 14572 4723
rect 14538 4515 14572 4531
rect 14326 4438 14342 4472
rect 14510 4438 14526 4472
rect 14166 4370 14200 4432
rect 14652 4370 14686 4432
rect 14166 4336 14262 4370
rect 14590 4336 14686 4370
rect 19636 4878 19732 4912
rect 20060 4878 20156 4912
rect 19636 4816 19670 4878
rect 20122 4816 20156 4878
rect 19796 4776 19812 4810
rect 19980 4776 19996 4810
rect 19750 4717 19784 4733
rect 19750 4525 19784 4541
rect 20008 4717 20042 4733
rect 20008 4525 20042 4541
rect 19796 4448 19812 4482
rect 19980 4448 19996 4482
rect 19636 4380 19670 4442
rect 20122 4380 20156 4442
rect 19636 4346 19732 4380
rect 20060 4346 20156 4380
rect 14166 3968 14262 4002
rect 14590 3968 14686 4002
rect 14166 3906 14200 3968
rect 14652 3906 14686 3968
rect 14326 3866 14342 3900
rect 14510 3866 14526 3900
rect 14280 3807 14314 3823
rect 14280 3615 14314 3631
rect 14538 3807 14572 3823
rect 14538 3615 14572 3631
rect 14326 3538 14342 3572
rect 14510 3538 14526 3572
rect 14166 3470 14200 3532
rect 14652 3470 14686 3532
rect 14166 3436 14262 3470
rect 14590 3436 14686 3470
rect 19636 3968 19732 4002
rect 20060 3968 20156 4002
rect 19636 3906 19670 3968
rect 20122 3906 20156 3968
rect 19796 3866 19812 3900
rect 19980 3866 19996 3900
rect 19750 3807 19784 3823
rect 19750 3615 19784 3631
rect 20008 3807 20042 3823
rect 20008 3615 20042 3631
rect 19796 3538 19812 3572
rect 19980 3538 19996 3572
rect 19636 3470 19670 3532
rect 20122 3470 20156 3532
rect 19636 3436 19732 3470
rect 20060 3436 20156 3470
rect 15366 3110 15462 3144
rect 15790 3110 15886 3144
rect 15366 3048 15400 3110
rect 15852 3048 15886 3110
rect 15526 3008 15542 3042
rect 15710 3008 15726 3042
rect 15480 2958 15514 2974
rect 15480 2766 15514 2782
rect 15738 2958 15772 2974
rect 15738 2766 15772 2782
rect 15526 2698 15542 2732
rect 15710 2698 15726 2732
rect 15366 2630 15400 2692
rect 15852 2630 15886 2692
rect 15366 2596 15462 2630
rect 15790 2596 15886 2630
rect 21446 3110 21542 3144
rect 21870 3110 21966 3144
rect 21446 3048 21480 3110
rect 21932 3048 21966 3110
rect 21606 3008 21622 3042
rect 21790 3008 21806 3042
rect 21560 2958 21594 2974
rect 21560 2766 21594 2782
rect 21818 2958 21852 2974
rect 21818 2766 21852 2782
rect 21606 2698 21622 2732
rect 21790 2698 21806 2732
rect 21446 2630 21480 2692
rect 21932 2630 21966 2692
rect 21446 2596 21542 2630
rect 21870 2596 21966 2630
rect 14426 2230 14522 2264
rect 14850 2230 14946 2264
rect 14426 2168 14460 2230
rect 14912 2168 14946 2230
rect 14586 2128 14602 2162
rect 14770 2128 14786 2162
rect 14540 2078 14574 2094
rect 14540 1886 14574 1902
rect 14798 2078 14832 2094
rect 14798 1886 14832 1902
rect 14586 1818 14602 1852
rect 14770 1818 14786 1852
rect 14426 1750 14460 1812
rect 14912 1750 14946 1812
rect 14426 1716 14522 1750
rect 14850 1716 14946 1750
rect 21456 2230 21552 2264
rect 21880 2230 21976 2264
rect 21456 2168 21490 2230
rect 21942 2168 21976 2230
rect 21616 2128 21632 2162
rect 21800 2128 21816 2162
rect 21570 2078 21604 2094
rect 21570 1886 21604 1902
rect 21828 2078 21862 2094
rect 21828 1886 21862 1902
rect 21616 1818 21632 1852
rect 21800 1818 21816 1852
rect 21456 1750 21490 1812
rect 21942 1750 21976 1812
rect 21456 1716 21552 1750
rect 21880 1716 21976 1750
rect 15814 1490 15830 1630
rect 16020 1490 16036 1630
<< viali >>
rect 15830 1490 16020 1630
<< metal1 >>
rect 15160 4780 19150 4830
rect 15110 4700 16935 4730
rect 15110 4240 15150 4700
rect 16610 4590 16690 4600
rect 16610 4580 16620 4590
rect 15380 4550 16620 4580
rect 16610 4520 16620 4550
rect 16680 4520 16690 4590
rect 16610 4510 16690 4520
rect 16980 4240 17020 4720
rect 17280 4410 17330 4780
rect 18110 4700 19380 4730
rect 17620 4590 17700 4600
rect 17620 4520 17630 4590
rect 17690 4580 17700 4590
rect 17690 4550 19110 4580
rect 17690 4520 17700 4550
rect 17620 4510 17700 4520
rect 17280 4400 17360 4410
rect 17280 4340 17290 4400
rect 17350 4340 17360 4400
rect 17280 4330 17360 4340
rect 17280 4300 17330 4330
rect 19260 4240 19380 4700
rect 13875 4110 19380 4240
rect 15110 3830 15150 4110
rect 15110 3800 16935 3830
rect 16610 3710 16710 3720
rect 16610 3680 16620 3710
rect 15380 3650 16620 3680
rect 16610 3620 16620 3650
rect 16700 3620 16710 3710
rect 16610 3610 16710 3620
rect 16980 3610 17020 4110
rect 19260 3830 19380 4110
rect 17280 3570 17310 3820
rect 18120 3800 19380 3830
rect 19260 3760 19380 3800
rect 17580 3710 17680 3720
rect 17580 3620 17590 3710
rect 17670 3680 17680 3710
rect 17670 3650 18940 3680
rect 17670 3620 17680 3650
rect 17580 3610 17680 3620
rect 15170 3520 19140 3570
rect 17280 3385 17310 3520
rect 17280 3355 17635 3385
rect 13880 3230 13990 3270
rect 13880 3190 15660 3230
rect 17605 3210 17635 3355
rect 13880 3160 13990 3190
rect 15620 2730 15660 3190
rect 16060 3170 21270 3210
rect 16060 2880 16100 3170
rect 16320 3080 16880 3120
rect 16170 2730 16180 2770
rect 15620 2700 16180 2730
rect 16270 2700 16280 2770
rect 15620 2690 16280 2700
rect 16320 2660 16360 3080
rect 16680 3040 16790 3050
rect 16680 2960 16690 3040
rect 16780 2960 16790 3040
rect 16680 2950 16790 2960
rect 15650 2620 16360 2660
rect 13880 2340 13990 2380
rect 13880 2300 15160 2340
rect 13880 2270 13990 2300
rect 15120 2160 15160 2300
rect 15120 2120 15620 2160
rect 15120 1920 15160 2120
rect 15380 1680 15420 2040
rect 15650 1900 15690 2620
rect 16575 2575 16625 2905
rect 16840 2660 16880 3080
rect 17100 2890 17140 3170
rect 17360 3080 17920 3120
rect 16920 2770 17030 2780
rect 16920 2700 16930 2770
rect 17020 2700 17030 2770
rect 16920 2690 17030 2700
rect 17180 2770 17300 2780
rect 17180 2700 17190 2770
rect 17290 2700 17300 2770
rect 17180 2690 17300 2700
rect 17360 2660 17400 3080
rect 17450 3040 17560 3050
rect 17450 2960 17460 3040
rect 17550 2960 17560 3040
rect 17450 2950 17560 2960
rect 17710 3040 17820 3050
rect 17710 2960 17720 3040
rect 17810 2960 17820 3040
rect 17710 2950 17820 2960
rect 16840 2620 17400 2660
rect 17605 2590 17655 2905
rect 17880 2660 17920 3080
rect 18130 2890 18170 3170
rect 18390 3080 18940 3120
rect 17950 2770 18070 2780
rect 17950 2700 17960 2770
rect 18060 2700 18070 2770
rect 17950 2690 18070 2700
rect 18220 2770 18340 2780
rect 18220 2700 18230 2770
rect 18330 2700 18340 2770
rect 18220 2690 18340 2700
rect 18390 2660 18430 3080
rect 18480 3040 18590 3050
rect 18480 2960 18490 3040
rect 18580 2960 18590 3040
rect 18480 2950 18590 2960
rect 18740 3040 18850 3050
rect 18740 2960 18750 3040
rect 18840 2960 18850 3040
rect 18740 2950 18850 2960
rect 17880 2620 18430 2660
rect 17570 2575 17655 2590
rect 18645 2575 18695 2945
rect 18900 2660 18940 3080
rect 19160 2890 19200 3170
rect 19420 3080 19980 3120
rect 18980 2770 19100 2780
rect 18980 2700 18990 2770
rect 19090 2700 19100 2770
rect 18980 2690 19100 2700
rect 19250 2770 19370 2780
rect 19250 2700 19260 2770
rect 19360 2700 19370 2770
rect 19250 2690 19370 2700
rect 19420 2660 19460 3080
rect 19520 3030 19630 3040
rect 19520 2950 19530 3030
rect 19620 2950 19630 3030
rect 19520 2940 19630 2950
rect 19770 3030 19880 3040
rect 19770 2950 19780 3030
rect 19870 2950 19880 3030
rect 19770 2940 19880 2950
rect 18900 2620 19460 2660
rect 19675 2575 19725 2905
rect 19940 2660 19980 3080
rect 20200 2890 20240 3170
rect 20450 3080 21010 3120
rect 20020 2770 20140 2780
rect 20020 2700 20030 2770
rect 20130 2700 20140 2770
rect 20020 2690 20140 2700
rect 20270 2770 20390 2780
rect 20270 2700 20280 2770
rect 20380 2700 20390 2770
rect 20270 2690 20390 2700
rect 20450 2660 20490 3080
rect 20540 3030 20650 3040
rect 20540 2950 20550 3030
rect 20640 2950 20650 3030
rect 20540 2940 20650 2950
rect 19940 2620 20490 2660
rect 20705 2575 20755 2905
rect 20970 2880 21010 3080
rect 21230 2900 21270 3170
rect 21050 2760 21170 2770
rect 16570 2560 20755 2575
rect 16570 2525 17270 2560
rect 17260 2480 17270 2525
rect 17370 2525 20755 2560
rect 20840 2530 20880 2730
rect 21050 2690 21060 2760
rect 21160 2690 21170 2760
rect 21050 2680 21170 2690
rect 17370 2480 17380 2525
rect 17570 2510 17650 2525
rect 20840 2490 21420 2530
rect 17100 2470 17200 2480
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 21380 2340 21420 2490
rect 16840 2300 22120 2340
rect 16060 2210 16620 2250
rect 16060 1680 16100 2210
rect 16130 1850 16180 1860
rect 16320 1850 16360 2080
rect 16130 1820 16360 1850
rect 16150 1810 16360 1820
rect 15380 1640 16100 1680
rect 16320 1680 16360 1810
rect 16580 1780 16620 2210
rect 16840 1950 16880 2300
rect 17100 2210 17660 2250
rect 17100 1780 17140 2210
rect 16580 1740 17140 1780
rect 17100 1708 17200 1710
rect 17100 1680 17113 1708
rect 16320 1640 17113 1680
rect 15710 1630 16100 1640
rect 15710 1490 15830 1630
rect 16020 1490 16100 1630
rect 17100 1633 17113 1640
rect 17188 1680 17200 1708
rect 17360 1680 17400 1960
rect 17620 1780 17660 2210
rect 17870 1970 17910 2300
rect 18130 2210 18690 2250
rect 18130 1780 18170 2210
rect 17620 1740 18170 1780
rect 18390 1680 18430 1970
rect 18650 1770 18690 2210
rect 18900 1950 18940 2300
rect 19160 2210 19720 2250
rect 19160 1770 19200 2210
rect 18650 1730 19200 1770
rect 19420 1680 19460 1960
rect 19680 1780 19720 2210
rect 19940 1960 19980 2300
rect 20190 2210 20750 2250
rect 20190 1780 20230 2210
rect 19680 1740 20230 1780
rect 20450 1680 20490 1960
rect 20710 1780 20750 2210
rect 20970 1950 21010 2300
rect 22010 2230 22120 2300
rect 21230 1780 21270 2000
rect 20710 1740 21270 1780
rect 17188 1640 20490 1680
rect 17188 1633 17200 1640
rect 17100 1620 17200 1633
rect 15710 1430 16100 1490
<< via1 >>
rect 16620 4520 16680 4590
rect 17630 4520 17690 4590
rect 17290 4340 17350 4400
rect 16620 3620 16700 3710
rect 17590 3620 17670 3710
rect 16180 2700 16270 2770
rect 16690 2960 16780 3040
rect 16930 2700 17020 2770
rect 17190 2700 17290 2770
rect 17460 2960 17550 3040
rect 17720 2960 17810 3040
rect 17960 2700 18060 2770
rect 18230 2700 18330 2770
rect 18490 2960 18580 3040
rect 18750 2960 18840 3040
rect 18990 2700 19090 2770
rect 19260 2700 19360 2770
rect 19530 2950 19620 3030
rect 19780 2950 19870 3030
rect 20030 2700 20130 2770
rect 20280 2700 20380 2770
rect 20550 2950 20640 3030
rect 17270 2480 17370 2560
rect 21060 2690 21160 2760
rect 17110 2390 17190 2470
rect 17113 1633 17188 1708
<< metal2 >>
rect 16610 4590 16690 4600
rect 16610 4520 16620 4590
rect 16680 4520 16690 4590
rect 16610 4510 16690 4520
rect 17620 4590 17700 4600
rect 17620 4520 17630 4590
rect 17690 4520 17700 4590
rect 17620 4510 17700 4520
rect 17280 4400 17360 4410
rect 17280 4340 17290 4400
rect 17350 4340 17360 4400
rect 16610 3710 16710 3720
rect 16610 3620 16620 3710
rect 16700 3620 16710 3710
rect 16610 3460 16710 3620
rect 16610 3360 16780 3460
rect 16680 3050 16780 3360
rect 17280 3330 17360 4340
rect 17405 3710 17680 3720
rect 17405 3620 17590 3710
rect 17670 3620 17680 3710
rect 17405 3610 17680 3620
rect 17270 3320 17370 3330
rect 17270 3230 17370 3240
rect 17405 3050 17515 3610
rect 16680 3040 17560 3050
rect 16680 2960 16690 3040
rect 16780 2960 17460 3040
rect 17550 2960 17560 3040
rect 16680 2950 17560 2960
rect 17710 3040 18590 3050
rect 17710 2960 17720 3040
rect 17810 2960 18490 3040
rect 18580 2960 18590 3040
rect 17710 2950 18590 2960
rect 18740 3040 19630 3050
rect 18740 2960 18750 3040
rect 18840 3030 19630 3040
rect 18840 2960 19530 3030
rect 18740 2950 19530 2960
rect 19620 2950 19630 3030
rect 18740 2940 19630 2950
rect 19770 3030 20650 3040
rect 19770 2950 19780 3030
rect 19870 2950 20550 3030
rect 20640 2950 20650 3030
rect 19770 2940 19880 2950
rect 20540 2940 20650 2950
rect 16180 2770 16270 2780
rect 16170 2700 16180 2760
rect 16920 2770 17030 2780
rect 16270 2740 16280 2760
rect 16920 2740 16930 2770
rect 16270 2700 16930 2740
rect 17020 2740 17030 2770
rect 17180 2770 17300 2780
rect 17020 2700 17040 2740
rect 16170 2690 17040 2700
rect 17180 2700 17190 2770
rect 17290 2700 17300 2770
rect 17180 2690 17300 2700
rect 17950 2770 18070 2780
rect 17950 2700 17960 2770
rect 18060 2700 18070 2770
rect 17950 2690 18070 2700
rect 18220 2770 19100 2780
rect 18220 2700 18230 2770
rect 18330 2700 18990 2770
rect 19090 2700 19100 2770
rect 18220 2690 19100 2700
rect 19250 2770 20140 2780
rect 19250 2700 19260 2770
rect 19360 2700 20030 2770
rect 20130 2700 20140 2770
rect 19250 2690 20140 2700
rect 20270 2770 21150 2780
rect 20270 2700 20280 2770
rect 20380 2760 21170 2770
rect 20380 2700 21060 2760
rect 20270 2690 21060 2700
rect 21160 2690 21170 2760
rect 21050 2680 21170 2690
rect 17260 2560 17380 2570
rect 17260 2480 17270 2560
rect 17370 2480 17380 2560
rect 17100 2470 17200 2480
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 17113 1710 17188 1718
rect 17100 1708 17200 1710
rect 17100 1633 17113 1708
rect 17188 1633 17200 1708
rect 17100 1620 17200 1633
<< via2 >>
rect 16620 4520 16680 4590
rect 17630 4520 17690 4590
rect 17270 3240 17370 3320
rect 17190 2700 17290 2770
rect 17960 2700 18060 2770
rect 17270 2480 17370 2560
rect 17110 2390 17190 2470
rect 17113 1633 17188 1708
<< metal3 >>
rect 16610 4590 17700 4600
rect 16610 4520 16620 4590
rect 16680 4520 17630 4590
rect 17690 4520 17700 4590
rect 16610 4510 17700 4520
rect 17110 3610 17190 4510
rect 17113 3390 17188 3610
rect 17100 3310 17110 3390
rect 17190 3310 17200 3390
rect 17260 3320 17380 3330
rect 17260 3240 17270 3320
rect 17370 3240 17380 3320
rect 17260 3230 17380 3240
rect 17180 2770 18070 2780
rect 17180 2700 17190 2770
rect 17290 2700 17960 2770
rect 18060 2700 18070 2770
rect 17180 2680 18070 2700
rect 17260 2560 17380 2570
rect 17113 2480 17188 2500
rect 17260 2480 17270 2560
rect 17370 2480 17380 2560
rect 17100 2470 17200 2480
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
rect 17113 1713 17188 2380
rect 17103 1710 17198 1713
rect 17100 1708 17200 1710
rect 17100 1633 17113 1708
rect 17188 1633 17200 1708
rect 17100 1620 17200 1633
<< via3 >>
rect 17110 3310 17190 3390
rect 17270 3240 17370 3320
rect 17270 2480 17370 2560
rect 17110 2390 17190 2470
<< metal4 >>
rect 17101 3390 17199 3399
rect 17100 3310 17110 3390
rect 17190 3310 17200 3390
rect 17100 3300 17200 3310
rect 17260 3320 17380 3340
rect 17101 2520 17199 3300
rect 17260 3240 17270 3320
rect 17370 3240 17380 3320
rect 17260 2560 17380 3240
rect 17100 2470 17200 2520
rect 17260 2480 17270 2560
rect 17370 2480 17380 2560
rect 17260 2470 17380 2480
rect 17100 2390 17110 2470
rect 17190 2390 17200 2470
rect 17100 2380 17200 2390
<< comment >>
rect 15530 4550 15940 4700
rect 17080 4540 17220 4700
rect 18220 4560 18630 4710
rect 15490 3640 15900 3790
rect 17100 3620 17240 3780
rect 18400 3630 18810 3780
rect 17940 2800 18620 2940
rect 15150 1910 15640 2070
rect 17940 1920 18620 2060
use sky130_fd_pr__nfet_01v8_CL66SD  sky130_fd_pr__nfet_01v8_CL66SD_0
timestamp 1661536226
transform 1 0 18667 0 1 2870
box -2747 -310 2747 310
use sky130_fd_pr__nfet_01v8_CL66SD  sky130_fd_pr__nfet_01v8_CL66SD_1
timestamp 1661536226
transform 1 0 18667 0 1 1990
box -2747 -310 2747 310
use sky130_fd_pr__nfet_01v8_GVTB53  sky130_fd_pr__nfet_01v8_GVTB53_0
timestamp 1661301161
transform 1 0 15405 0 1 1990
box -425 -310 425 310
use sky130_fd_pr__pfet_01v8_8C4HA7  sky130_fd_pr__pfet_01v8_8C4HA7_0
timestamp 1661301161
transform 1 0 15792 0 1 3719
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_8L4H97  sky130_fd_pr__pfet_01v8_8L4H97_0
timestamp 1661301161
transform 1 0 15792 0 1 4619
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_8LYGA7  sky130_fd_pr__pfet_01v8_8LYGA7_0
timestamp 1661301161
transform -1 0 18532 0 1 4619
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_8LYGA7  sky130_fd_pr__pfet_01v8_8LYGA7_1
timestamp 1661301161
transform -1 0 18532 0 1 3719
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_BLSBYX  sky130_fd_pr__pfet_01v8_BLSBYX_0
timestamp 1661301161
transform 1 0 17156 0 1 4619
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_BLSBYX  sky130_fd_pr__pfet_01v8_BLSBYX_1
timestamp 1661301161
transform 1 0 17156 0 1 3719
box -296 -319 296 319
<< labels >>
flabel metal1 19710 1650 19750 1660 0 FreeSans 800 0 0 0 net1
flabel metal1 15710 1490 15820 1600 0 FreeSans 1600 0 0 0 gnd
port 4 nsew
flabel comment 15220 1920 15340 2050 0 FreeSans 800 0 0 0 M10
flabel comment 15470 1920 15590 2050 0 FreeSans 800 0 0 0 M5
flabel comment 15490 3640 15900 3790 0 FreeSans 800 0 0 0 M6_1
flabel comment 18220 4560 18630 4710 0 FreeSans 800 0 0 0 M8_2
flabel comment 15530 4550 15940 4700 0 FreeSans 800 0 0 0 M8_1
flabel comment 17080 4540 17220 4700 0 FreeSans 800 0 0 0 M3
flabel comment 18400 3630 18810 3780 0 FreeSans 800 0 0 0 M6_2
flabel metal2 17320 4070 17320 4070 0 FreeSans 800 0 0 0 net2
flabel comment 17100 3620 17240 3780 0 FreeSans 800 0 0 0 M4
flabel metal1 15670 2390 15680 2410 0 FreeSans 800 0 0 0 net4
flabel comment 17940 1920 18620 2060 0 FreeSans 800 0 0 0 M9_M7
flabel comment 17940 2800 18620 2940 0 FreeSans 800 0 0 0 M1_M2
flabel metal1 17600 3360 17620 3380 0 FreeSans 800 0 0 0 net3
flabel metal1 13880 4120 13990 4230 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 13880 3160 13990 3270 0 FreeSans 1600 0 0 0 in
port 3 nsew
flabel metal1 13880 2270 13990 2380 0 FreeSans 1600 0 0 0 ib
port 1 nsew
flabel metal1 22010 2230 22120 2340 0 FreeSans 1600 0 0 0 out
port 2 nsew
<< end >>
