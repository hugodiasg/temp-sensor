magic
tech sky130A
magscale 1 2
timestamp 1645645281
<< metal4 >>
rect -2629 7709 2629 7750
rect -2629 2691 2373 7709
rect 2609 2691 2629 7709
rect -2629 2650 2629 2691
rect -2629 2509 2629 2550
rect -2629 -2509 2373 2509
rect 2609 -2509 2629 2509
rect -2629 -2550 2629 -2509
rect -2629 -2691 2629 -2650
rect -2629 -7709 2373 -2691
rect 2609 -7709 2629 -2691
rect -2629 -7750 2629 -7709
<< via4 >>
rect 2373 2691 2609 7709
rect 2373 -2509 2609 2509
rect 2373 -7709 2609 -2691
<< mimcap2 >>
rect -2529 7610 2371 7650
rect -2529 2790 -2007 7610
rect 1849 2790 2371 7610
rect -2529 2750 2371 2790
rect -2529 2410 2371 2450
rect -2529 -2410 -2007 2410
rect 1849 -2410 2371 2410
rect -2529 -2450 2371 -2410
rect -2529 -2790 2371 -2750
rect -2529 -7610 -2007 -2790
rect 1849 -7610 2371 -2790
rect -2529 -7650 2371 -7610
<< mimcap2contact >>
rect -2007 2790 1849 7610
rect -2007 -2410 1849 2410
rect -2007 -7610 1849 -2790
<< metal5 >>
rect -239 7634 81 7800
rect 2331 7709 2651 7800
rect -2031 7610 1873 7634
rect -2031 2790 -2007 7610
rect 1849 2790 1873 7610
rect -2031 2766 1873 2790
rect -239 2434 81 2766
rect 2331 2691 2373 7709
rect 2609 2691 2651 7709
rect 2331 2509 2651 2691
rect -2031 2410 1873 2434
rect -2031 -2410 -2007 2410
rect 1849 -2410 1873 2410
rect -2031 -2434 1873 -2410
rect -239 -2766 81 -2434
rect 2331 -2509 2373 2509
rect 2609 -2509 2651 2509
rect 2331 -2691 2651 -2509
rect -2031 -2790 1873 -2766
rect -2031 -7610 -2007 -2790
rect 1849 -7610 1873 -2790
rect -2031 -7634 1873 -7610
rect -239 -7800 81 -7634
rect 2331 -7709 2373 -2691
rect 2609 -7709 2651 -2691
rect 2331 -7800 2651 -7709
<< properties >>
string FIXED_BBOX -2629 2650 2471 7750
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.5 l 24.5 val 1.219k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
