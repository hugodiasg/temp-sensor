magic
tech sky130A
magscale 1 2
timestamp 1656877262
<< mvpsubdiff >>
rect 6561 -7206 6585 -7006
rect 6945 -7206 6969 -7006
<< mvpsubdiffcont >>
rect 6585 -7206 6945 -7006
<< locali >>
rect 6569 -7206 6585 -7006
rect 6945 -7206 6961 -7006
<< viali >>
rect 6585 -7206 6945 -7006
<< metal1 >>
rect 6300 16620 9480 16640
rect 6300 16140 8840 16620
rect 9460 16140 9480 16620
rect 6300 16120 9480 16140
rect 7700 -1680 9360 -1640
rect 7700 -2760 7720 -1680
rect 8600 -2180 9360 -1680
rect 10360 -1660 11560 -1620
rect 10360 -2100 10960 -1660
rect 11540 -2100 11560 -1660
rect 10360 -2158 11560 -2100
rect 10360 -2160 10954 -2158
rect 8600 -2760 8680 -2180
rect 8860 -2580 10360 -2240
rect 7700 -2800 8680 -2760
rect 9960 -2800 10360 -2580
rect 6340 -4480 9760 -2800
rect 9880 -3360 10360 -2800
rect 9880 -3740 10660 -3360
rect 9880 -4480 10360 -3740
rect 9718 -4646 9884 -4572
rect 9720 -5160 9880 -4646
rect 6340 -5360 9880 -5160
rect 10480 -6765 10660 -3740
rect 6573 -7006 6957 -7000
rect 10480 -7006 10664 -6765
rect 6345 -7206 6585 -7006
rect 6945 -7206 10664 -7006
rect 6573 -7212 6957 -7206
<< via1 >>
rect 8840 16140 9460 16620
rect 7720 -2760 8600 -1680
rect 10960 -2100 11540 -1660
<< metal2 >>
rect 8820 16620 9480 16640
rect 8820 16140 8840 16620
rect 9460 16140 9480 16620
rect 8820 16120 9480 16140
rect 7700 -1640 8600 -1620
rect 7700 -1680 8660 -1640
rect 7700 -2760 7720 -1680
rect 8600 -2760 8660 -1680
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
rect 7700 -2820 8660 -2760
<< via2 >>
rect 8840 16140 9460 16620
rect 7720 -2760 8600 -1680
rect 10960 -2100 11540 -1660
<< metal3 >>
rect 8820 16620 9480 16640
rect 8820 16140 8840 16620
rect 9460 16140 9480 16620
rect 8820 16120 9480 16140
rect 7700 -1640 8600 -1620
rect 7700 -1680 8660 -1640
rect 7700 -2760 7720 -1680
rect 8600 -2760 8660 -1680
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
rect 7700 -2820 8660 -2760
<< via3 >>
rect 8840 16140 9460 16620
rect 7720 -2760 8600 -1680
rect 10960 -2100 11540 -1660
<< metal4 >>
rect 8820 16620 9480 16640
rect 8820 16140 8840 16620
rect 9460 16140 9480 16620
rect 8820 16120 9480 16140
rect 7020 9040 12260 9420
rect 7020 3840 12260 4260
rect 7700 -1640 8600 -329
rect 9220 -380 15380 1980
rect 7700 -1680 8660 -1640
rect 7700 -2760 7720 -1680
rect 8600 -2760 8660 -1680
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
rect 7700 -2820 8660 -2760
rect 13020 -6420 15380 -380
rect 13020 -8780 30458 -6420
<< via4 >>
rect 8840 16140 9460 16620
rect 10960 -2100 11540 -1660
<< metal5 >>
rect 8819 17560 12940 17562
rect 13860 17560 15123 17562
rect 8819 16644 15123 17560
rect 8816 16620 15123 16644
rect 8816 16140 8840 16620
rect 9460 16140 15123 16620
rect 8816 16116 15123 16140
rect 8819 15200 15123 16116
rect 8819 12219 11181 15200
rect 9200 12200 10400 12219
rect 10940 -1600 11580 -338
rect 10920 -1660 11580 -1600
rect 10920 -2100 10960 -1660
rect 11540 -2100 11580 -1660
rect 10920 -2140 11580 -2100
use l0_0  l0_0_0
timestamp 1647142466
transform 1 0 -24400 0 1 -45638
box 39200 36838 63200 63200
use sky130_fd_pr__cap_mim_m3_2_97K3D8  sky130_fd_pr__cap_mim_m3_2_97K3D8_0
timestamp 1647142466
transform -1 0 9641 0 1 6632
box -2619 -7770 2641 7770
use sky130_fd_pr__nfet_g5v0d10v5_PWYS4E  sky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0
timestamp 1647142466
transform 1 0 9796 0 1 -3646
box -278 -1128 278 1128
use sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN  sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0
timestamp 1647142466
transform 0 1 9872 -1 0 -2093
box -201 -1098 201 1098
<< labels >>
flabel metal1 6340 -3040 6540 -2840 0 FreeSans 9600 0 0 0 out
port 2 nsew
flabel metal1 6340 -5360 6540 -5160 0 FreeSans 9600 0 0 0 in
port 1 nsew
flabel metal1 6340 16440 6540 16640 0 FreeSans 9600 0 0 0 vd
port 3 nsew
flabel metal1 6345 -7206 6545 -7006 0 FreeSans 9600 0 0 0 gnd
port 0 nsew
<< end >>
