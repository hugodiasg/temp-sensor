** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sch
.subckt ask-modulator gnd in out vd
*.PININFO gnd:B in:I out:O vd:B
XM2 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 vd out sky130_fd_pr__cap_mim_m3_2 W=24.5 L=24.5 MF=1 m=1
XC2 vd out sky130_fd_pr__cap_mim_m3_2 W=24.5 L=24.5 MF=1 m=1
XC3 vd out sky130_fd_pr__cap_mim_m3_2 W=24.5 L=24.5 MF=1 m=1
XR1 out vd gnd sky130_fd_pr__res_high_po_5p73 L=0.5 mult=1 m=1
L1 vd out 1n m=1
**** begin user architecture code



**** end user architecture code
.ends
.end
