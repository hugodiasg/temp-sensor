magic
tech sky130A
magscale 1 2
timestamp 1700007007
<< nwell >>
rect -1457 -319 1457 319
<< pmos >>
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
<< pdiff >>
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
<< pdiffc >>
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
<< nsubdiff >>
rect -1421 249 -1325 283
rect 1325 249 1421 283
rect -1421 187 -1387 249
rect 1387 187 1421 249
rect -1421 -249 -1387 -187
rect 1387 -249 1421 -187
rect -1421 -283 -1325 -249
rect 1325 -283 1421 -249
<< nsubdiffcont >>
rect -1325 249 1325 283
rect -1421 -187 -1387 187
rect 1387 -187 1421 187
rect -1325 -283 1325 -249
<< poly >>
rect -1261 181 -1061 197
rect -1261 147 -1245 181
rect -1077 147 -1061 181
rect -1261 100 -1061 147
rect -1003 181 -803 197
rect -1003 147 -987 181
rect -819 147 -803 181
rect -1003 100 -803 147
rect -745 181 -545 197
rect -745 147 -729 181
rect -561 147 -545 181
rect -745 100 -545 147
rect -487 181 -287 197
rect -487 147 -471 181
rect -303 147 -287 181
rect -487 100 -287 147
rect -229 181 -29 197
rect -229 147 -213 181
rect -45 147 -29 181
rect -229 100 -29 147
rect 29 181 229 197
rect 29 147 45 181
rect 213 147 229 181
rect 29 100 229 147
rect 287 181 487 197
rect 287 147 303 181
rect 471 147 487 181
rect 287 100 487 147
rect 545 181 745 197
rect 545 147 561 181
rect 729 147 745 181
rect 545 100 745 147
rect 803 181 1003 197
rect 803 147 819 181
rect 987 147 1003 181
rect 803 100 1003 147
rect 1061 181 1261 197
rect 1061 147 1077 181
rect 1245 147 1261 181
rect 1061 100 1261 147
rect -1261 -147 -1061 -100
rect -1261 -181 -1245 -147
rect -1077 -181 -1061 -147
rect -1261 -197 -1061 -181
rect -1003 -147 -803 -100
rect -1003 -181 -987 -147
rect -819 -181 -803 -147
rect -1003 -197 -803 -181
rect -745 -147 -545 -100
rect -745 -181 -729 -147
rect -561 -181 -545 -147
rect -745 -197 -545 -181
rect -487 -147 -287 -100
rect -487 -181 -471 -147
rect -303 -181 -287 -147
rect -487 -197 -287 -181
rect -229 -147 -29 -100
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect -229 -197 -29 -181
rect 29 -147 229 -100
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 29 -197 229 -181
rect 287 -147 487 -100
rect 287 -181 303 -147
rect 471 -181 487 -147
rect 287 -197 487 -181
rect 545 -147 745 -100
rect 545 -181 561 -147
rect 729 -181 745 -147
rect 545 -197 745 -181
rect 803 -147 1003 -100
rect 803 -181 819 -147
rect 987 -181 1003 -147
rect 803 -197 1003 -181
rect 1061 -147 1261 -100
rect 1061 -181 1077 -147
rect 1245 -181 1261 -147
rect 1061 -197 1261 -181
<< polycont >>
rect -1245 147 -1077 181
rect -987 147 -819 181
rect -729 147 -561 181
rect -471 147 -303 181
rect -213 147 -45 181
rect 45 147 213 181
rect 303 147 471 181
rect 561 147 729 181
rect 819 147 987 181
rect 1077 147 1245 181
rect -1245 -181 -1077 -147
rect -987 -181 -819 -147
rect -729 -181 -561 -147
rect -471 -181 -303 -147
rect -213 -181 -45 -147
rect 45 -181 213 -147
rect 303 -181 471 -147
rect 561 -181 729 -147
rect 819 -181 987 -147
rect 1077 -181 1245 -147
<< locali >>
rect -1421 249 -1325 283
rect 1325 249 1421 283
rect -1421 187 -1387 249
rect 1387 187 1421 249
rect -1261 147 -1245 181
rect -1077 147 -1061 181
rect -1003 147 -987 181
rect -819 147 -803 181
rect -745 147 -729 181
rect -561 147 -545 181
rect -487 147 -471 181
rect -303 147 -287 181
rect -229 147 -213 181
rect -45 147 -29 181
rect 29 147 45 181
rect 213 147 229 181
rect 287 147 303 181
rect 471 147 487 181
rect 545 147 561 181
rect 729 147 745 181
rect 803 147 819 181
rect 987 147 1003 181
rect 1061 147 1077 181
rect 1245 147 1261 181
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect -1261 -181 -1245 -147
rect -1077 -181 -1061 -147
rect -1003 -181 -987 -147
rect -819 -181 -803 -147
rect -745 -181 -729 -147
rect -561 -181 -545 -147
rect -487 -181 -471 -147
rect -303 -181 -287 -147
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 287 -181 303 -147
rect 471 -181 487 -147
rect 545 -181 561 -147
rect 729 -181 745 -147
rect 803 -181 819 -147
rect 987 -181 1003 -147
rect 1061 -181 1077 -147
rect 1245 -181 1261 -147
rect -1421 -249 -1387 -187
rect 1387 -249 1421 -187
rect -1421 -283 -1325 -249
rect 1325 -283 1421 -249
<< viali >>
rect -1245 147 -1077 181
rect -987 147 -819 181
rect -729 147 -561 181
rect -471 147 -303 181
rect -213 147 -45 181
rect 45 147 213 181
rect 303 147 471 181
rect 561 147 729 181
rect 819 147 987 181
rect 1077 147 1245 181
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect -1245 -181 -1077 -147
rect -987 -181 -819 -147
rect -729 -181 -561 -147
rect -471 -181 -303 -147
rect -213 -181 -45 -147
rect 45 -181 213 -147
rect 303 -181 471 -147
rect 561 -181 729 -147
rect 819 -181 987 -147
rect 1077 -181 1245 -147
<< metal1 >>
rect -1257 181 -1065 187
rect -1257 147 -1245 181
rect -1077 147 -1065 181
rect -1257 141 -1065 147
rect -999 181 -807 187
rect -999 147 -987 181
rect -819 147 -807 181
rect -999 141 -807 147
rect -741 181 -549 187
rect -741 147 -729 181
rect -561 147 -549 181
rect -741 141 -549 147
rect -483 181 -291 187
rect -483 147 -471 181
rect -303 147 -291 181
rect -483 141 -291 147
rect -225 181 -33 187
rect -225 147 -213 181
rect -45 147 -33 181
rect -225 141 -33 147
rect 33 181 225 187
rect 33 147 45 181
rect 213 147 225 181
rect 33 141 225 147
rect 291 181 483 187
rect 291 147 303 181
rect 471 147 483 181
rect 291 141 483 147
rect 549 181 741 187
rect 549 147 561 181
rect 729 147 741 181
rect 549 141 741 147
rect 807 181 999 187
rect 807 147 819 181
rect 987 147 999 181
rect 807 141 999 147
rect 1065 181 1257 187
rect 1065 147 1077 181
rect 1245 147 1257 181
rect 1065 141 1257 147
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect -1257 -147 -1065 -141
rect -1257 -181 -1245 -147
rect -1077 -181 -1065 -147
rect -1257 -187 -1065 -181
rect -999 -147 -807 -141
rect -999 -181 -987 -147
rect -819 -181 -807 -147
rect -999 -187 -807 -181
rect -741 -147 -549 -141
rect -741 -181 -729 -147
rect -561 -181 -549 -147
rect -741 -187 -549 -181
rect -483 -147 -291 -141
rect -483 -181 -471 -147
rect -303 -181 -291 -147
rect -483 -187 -291 -181
rect -225 -147 -33 -141
rect -225 -181 -213 -147
rect -45 -181 -33 -147
rect -225 -187 -33 -181
rect 33 -147 225 -141
rect 33 -181 45 -147
rect 213 -181 225 -147
rect 33 -187 225 -181
rect 291 -147 483 -141
rect 291 -181 303 -147
rect 471 -181 483 -147
rect 291 -187 483 -181
rect 549 -147 741 -141
rect 549 -181 561 -147
rect 729 -181 741 -147
rect 549 -187 741 -181
rect 807 -147 999 -141
rect 807 -181 819 -147
rect 987 -181 999 -147
rect 807 -187 999 -181
rect 1065 -147 1257 -141
rect 1065 -181 1077 -147
rect 1245 -181 1257 -147
rect 1065 -187 1257 -181
<< properties >>
string FIXED_BBOX -1404 -266 1404 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
