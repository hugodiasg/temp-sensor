magic
tech sky130A
magscale 1 2
timestamp 1644600357
<< mvpsubdiff >>
rect 6760 -4260 6940 -4236
rect 6760 -4484 6940 -4460
<< mvpsubdiffcont >>
rect 6760 -4460 6940 -4260
<< viali >>
rect 6760 -4260 6940 -4240
rect 6760 -4460 6940 -4260
rect 6760 -4480 6940 -4460
<< metal1 >>
rect 2740 -1340 5760 -1240
rect 2740 -1700 2780 -1340
rect 3500 -1700 5760 -1340
rect 2740 -1780 5760 -1700
rect 6760 -1320 10400 -1220
rect 6760 -1680 9640 -1320
rect 10360 -1680 10400 -1320
rect 6760 -1760 10400 -1680
rect 4880 -2400 5080 -1780
rect 5260 -2180 6760 -1840
rect 6360 -2400 6760 -2180
rect 4880 -2920 6160 -2400
rect 4620 -3300 6160 -2920
rect 4620 -4520 4780 -3300
rect 4880 -4100 6160 -3300
rect 6280 -2960 6760 -2400
rect 6280 -3340 7060 -2960
rect 6280 -4100 6760 -3340
rect 6120 -4520 6280 -4140
rect 6900 -4220 7060 -3340
rect 6740 -4240 7060 -4220
rect 6740 -4480 6760 -4240
rect 6940 -4480 7060 -4240
rect 6740 -4500 7060 -4480
rect 7360 -4500 7520 -1760
rect 6740 -4520 7080 -4500
rect 4600 -4720 4800 -4520
rect 6100 -4720 6300 -4520
rect 6880 -4700 7080 -4520
rect 7340 -4700 7540 -4500
<< via1 >>
rect 2780 -1700 3500 -1340
rect 9640 -1680 10360 -1320
<< metal2 >>
rect 2740 -1340 3540 -1300
rect 2740 -1700 2780 -1340
rect 3500 -1700 3540 -1340
rect 2740 -1780 3540 -1700
rect 9600 -1320 10400 -1280
rect 9600 -1680 9640 -1320
rect 10360 -1680 10400 -1320
rect 9600 -1760 10400 -1680
<< via2 >>
rect 2780 -1700 3500 -1340
rect 9640 -1680 10360 -1320
<< metal3 >>
rect 2740 -1340 3540 -1300
rect 2740 -1700 2780 -1340
rect 3500 -1700 3540 -1340
rect 2740 -1780 3540 -1700
rect 9600 -1320 10400 -1280
rect 9600 -1680 9640 -1320
rect 10360 -1680 10400 -1320
rect 9600 -1760 10400 -1680
<< via3 >>
rect 2780 -1700 3500 -1340
rect 9640 -1680 10360 -1320
<< metal4 >>
rect 2740 15600 3540 15660
rect 2740 14800 17200 15600
rect 2740 -1340 3540 14800
rect 6000 13600 6800 14800
rect 2740 -1700 2780 -1340
rect 3500 -1700 3540 -1340
rect 2740 -1780 3540 -1700
rect 9600 -1320 10400 -1280
rect 9600 -1680 9640 -1320
rect 10360 -1680 10400 -1320
rect 9600 -1760 10400 -1680
<< via4 >>
rect 9640 -1680 10360 -1320
<< metal5 >>
rect 6120 13600 12200 14400
rect 9600 -1320 10400 13600
rect 9600 -1680 9640 -1320
rect 10360 -1680 10400 -1320
rect 9600 -1760 10400 -1680
use sky130_fd_pr__cap_mim_m3_2_QKF9RA  XC0
timestamp 1644600357
transform -1 0 6101 0 1 6950
box -2479 -7350 2501 7350
use sky130_fd_pr__res_xhigh_po_0p35_NVRUDW  XR1
timestamp 1644594744
transform 0 1 6258 -1 0 -1699
box -201 -1098 201 1098
use sky130_fd_pr__nfet_g5v0d10v5_ML7W5H  XM1
timestamp 1644594744
transform -1 0 6218 0 1 -3232
box -278 -1128 278 1128
use l0  x1
timestamp 1644598236
transform 1 0 10916 0 1 -1459
box -116 -141 15884 16659
<< labels >>
flabel metal1 6100 -4720 6300 -4520 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 4600 -4720 4800 -4520 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 6880 -4700 7080 -4500 0 FreeSans 128 0 0 0 gnd
port 0 nsew
flabel metal1 7340 -4700 7540 -4500 0 FreeSans 128 0 0 0 vd
port 3 nsew
<< end >>
