magic
tech sky130A
magscale 1 2
timestamp 1669420244
<< nwell >>
rect -256 -1419 256 1419
<< pmos >>
rect -60 -1200 60 1200
<< pdiff >>
rect -118 1188 -60 1200
rect -118 -1188 -106 1188
rect -72 -1188 -60 1188
rect -118 -1200 -60 -1188
rect 60 1188 118 1200
rect 60 -1188 72 1188
rect 106 -1188 118 1188
rect 60 -1200 118 -1188
<< pdiffc >>
rect -106 -1188 -72 1188
rect 72 -1188 106 1188
<< nsubdiff >>
rect -220 1349 -124 1383
rect 124 1349 220 1383
rect -220 1287 -186 1349
rect 186 1287 220 1349
rect -220 -1349 -186 -1287
rect 186 -1349 220 -1287
rect -220 -1383 -124 -1349
rect 124 -1383 220 -1349
<< nsubdiffcont >>
rect -124 1349 124 1383
rect -220 -1287 -186 1287
rect 186 -1287 220 1287
rect -124 -1383 124 -1349
<< poly >>
rect -60 1281 60 1297
rect -60 1247 -44 1281
rect 44 1247 60 1281
rect -60 1200 60 1247
rect -60 -1247 60 -1200
rect -60 -1281 -44 -1247
rect 44 -1281 60 -1247
rect -60 -1297 60 -1281
<< polycont >>
rect -44 1247 44 1281
rect -44 -1281 44 -1247
<< locali >>
rect -220 1349 -124 1383
rect 124 1349 220 1383
rect -220 1287 -186 1349
rect 186 1287 220 1349
rect -60 1247 -44 1281
rect 44 1247 60 1281
rect -106 1188 -72 1204
rect -106 -1204 -72 -1188
rect 72 1188 106 1204
rect 72 -1204 106 -1188
rect -60 -1281 -44 -1247
rect 44 -1281 60 -1247
rect -220 -1349 -186 -1287
rect 186 -1349 220 -1287
rect -220 -1383 -124 -1349
rect 124 -1383 220 -1349
<< viali >>
rect -44 1247 44 1281
rect -106 -1188 -72 1188
rect 72 -1188 106 1188
rect -44 -1281 44 -1247
<< metal1 >>
rect -56 1281 56 1287
rect -56 1247 -44 1281
rect 44 1247 56 1281
rect -56 1241 56 1247
rect -112 1188 -66 1200
rect -112 -1188 -106 1188
rect -72 -1188 -66 1188
rect -112 -1200 -66 -1188
rect 66 1188 112 1200
rect 66 -1188 72 1188
rect 106 -1188 112 1188
rect 66 -1200 112 -1188
rect -56 -1247 56 -1241
rect -56 -1281 -44 -1247
rect 44 -1281 56 -1247
rect -56 -1287 56 -1281
<< properties >>
string FIXED_BBOX -203 -1366 203 1366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 12 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
