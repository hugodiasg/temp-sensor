magic
tech sky130A
magscale 1 2
timestamp 1646426626
<< metal4 >>
rect -2614 7664 2614 7705
rect -2614 2676 2358 7664
rect 2594 2676 2614 7664
rect -2614 2635 2614 2676
rect -2614 2494 2614 2535
rect -2614 -2494 2358 2494
rect 2594 -2494 2614 2494
rect -2614 -2535 2614 -2494
rect -2614 -2676 2614 -2635
rect -2614 -7664 2358 -2676
rect 2594 -7664 2614 -2676
rect -2614 -7705 2614 -7664
<< via4 >>
rect 2358 2676 2594 7664
rect 2358 -2494 2594 2494
rect 2358 -7664 2594 -2676
<< mimcap2 >>
rect -2514 7565 2356 7605
rect -2514 2775 -1995 7565
rect 1837 2775 2356 7565
rect -2514 2735 2356 2775
rect -2514 2395 2356 2435
rect -2514 -2395 -1995 2395
rect 1837 -2395 2356 2395
rect -2514 -2435 2356 -2395
rect -2514 -2775 2356 -2735
rect -2514 -7565 -1995 -2775
rect 1837 -7565 2356 -2775
rect -2514 -7605 2356 -7565
<< mimcap2contact >>
rect -1995 2775 1837 7565
rect -1995 -2395 1837 2395
rect -1995 -7565 1837 -2775
<< metal5 >>
rect -239 7589 81 7755
rect 2316 7664 2636 7755
rect -2019 7565 1861 7589
rect -2019 2775 -1995 7565
rect 1837 2775 1861 7565
rect -2019 2751 1861 2775
rect -239 2419 81 2751
rect 2316 2676 2358 7664
rect 2594 2676 2636 7664
rect 2316 2494 2636 2676
rect -2019 2395 1861 2419
rect -2019 -2395 -1995 2395
rect 1837 -2395 1861 2395
rect -2019 -2419 1861 -2395
rect -239 -2751 81 -2419
rect 2316 -2494 2358 2494
rect 2594 -2494 2636 2494
rect 2316 -2676 2636 -2494
rect -2019 -2775 1861 -2751
rect -2019 -7565 -1995 -2775
rect 1837 -7565 1861 -2775
rect -2019 -7589 1861 -7565
rect -239 -7755 81 -7589
rect 2316 -7664 2358 -2676
rect 2594 -7664 2636 -2676
rect 2316 -7755 2636 -7664
<< properties >>
string FIXED_BBOX -2614 2635 2456 7705
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.35 l 24.35 val 1.204k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
