** sch_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/dff_tb-tran.sch
**.subckt dff_tb-tran
vclk clk GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 50ns 100ns)
VDD vd GND 1.8
vin in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 1.5us 3us)
x1 clk in vd GND GND VD VD q qn sky130_fd_sc_hd__dfrbp_1
**** begin user architecture code

*cmd step stop
.tran 0.5n 5u
.control
set color0=white
set color1=black
set temp=27
destroy all
run

plot in
plot clk
plot q qn


.endc

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
