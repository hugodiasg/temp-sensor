magic
tech sky130A
timestamp 1644950992
<< metal4 >>
rect -600 1479 1500 1500
rect -600 920 918 1479
rect 1481 920 1500 1479
rect -600 900 1500 920
<< via4 >>
rect 918 920 1481 1479
<< metal5 >>
rect 0 14400 15000 15000
rect 0 13500 14100 14100
rect 0 600 600 13500
rect 13500 1500 14100 13500
rect 900 1479 14100 1500
rect 900 920 918 1479
rect 1481 920 14100 1479
rect 900 900 14100 920
rect 14400 600 15000 14400
rect 0 0 15000 600
<< end >>
