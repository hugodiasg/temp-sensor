** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator_tb-tran.sch
**.subckt ask-modulator_tb-tran
Vdd vd GND 3.3
Vin in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 6ns 12ns)
x1 vd out in GND ask-modulator
**** begin user architecture code

.tran 0.01n 8n
.control
destroy all
run
let id =-i(vdd)
let z_rlc= (vd-out)/id
let z_nmos=out/id
let z_out=z_rlc*z_nmos/(z_rlc+z_nmos)
plot z_out
plot id
plot in
plot out
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  ask-modulator.sym # of pins=4
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sch
.subckt ask-modulator  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XM2 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=1 W=21 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
L0 vd out 5.097n m=1
XC0 vd out sky130_fd_pr__cap_mim_m3_1 W=19.75 L=19.75 MF=1 m=1
XR0 out vd gnd sky130_fd_pr__res_high_po_5p73 L=0.5 mult=1 m=1
.ends

.GLOBAL GND
.end
