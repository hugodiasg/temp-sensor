magic
tech sky130A
magscale 1 2
timestamp 1675974324
use sky130_fd_pr__cap_mim_m3_2_MVDWNN  XC0
timestamp 1675895675
transform 1 0 -8807 0 1 -7080
box -14145 -12600 14167 12600
use sky130_fd_pr__cap_mim_m3_2_M62EV7  XC1
timestamp 1675895675
transform 1 0 22130 0 1 -5826
box -15145 -13600 15167 13600
use l0  l0_0
timestamp 1675896714
transform 1 0 -44497 0 1 -81349
box 42526 43199 62561 59200
<< end >>
