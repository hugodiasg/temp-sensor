magic
tech sky130A
magscale 1 2
timestamp 1644161670
<< error_p >>
rect 2133 -7650 2429 7650
rect 2453 2821 2749 7601
rect 2453 2599 2773 2821
rect 2453 2279 2773 2501
rect 2453 -2279 2749 2279
rect 2453 -2501 2773 -2279
rect 2453 -2821 2773 -2599
rect 2453 -7601 2749 -2821
<< metal4 >>
rect -2751 7559 2751 7600
rect -2751 2641 2495 7559
rect 2731 2641 2751 7559
rect -2751 2600 2751 2641
rect -2751 2459 2751 2500
rect -2751 -2459 2495 2459
rect 2731 -2459 2751 2459
rect -2751 -2500 2751 -2459
rect -2751 -2641 2751 -2600
rect -2751 -7559 2495 -2641
rect 2731 -7559 2751 -2641
rect -2751 -7600 2751 -7559
<< via4 >>
rect 2495 2641 2731 7559
rect 2495 -2459 2731 2459
rect 2495 -7559 2731 -2641
<< mimcap2 >>
rect -2651 7460 2149 7500
rect -2651 2740 -2611 7460
rect 2109 2740 2149 7460
rect -2651 2700 2149 2740
rect -2651 2360 2149 2400
rect -2651 -2360 -2611 2360
rect 2109 -2360 2149 2360
rect -2651 -2400 2149 -2360
rect -2651 -2740 2149 -2700
rect -2651 -7460 -2611 -2740
rect 2109 -7460 2149 -2740
rect -2651 -7500 2149 -7460
<< mimcap2contact >>
rect -2611 2740 2109 7460
rect -2611 -2360 2109 2360
rect -2611 -7460 2109 -2740
<< metal5 >>
rect -411 7484 -91 7650
rect 2109 7484 2429 7650
rect -2635 7460 2429 7484
rect -2635 2740 -2611 7460
rect 2109 2740 2429 7460
rect -2635 2716 2429 2740
rect -411 2384 -91 2716
rect 2109 2384 2429 2716
rect 2453 7559 2773 7601
rect 2453 2641 2495 7559
rect 2731 2641 2773 7559
rect 2453 2599 2773 2641
rect -2635 2360 2429 2384
rect -2635 -2360 -2611 2360
rect 2109 -2360 2429 2360
rect -2635 -2384 2429 -2360
rect -411 -2716 -91 -2384
rect 2109 -2716 2429 -2384
rect 2453 2459 2773 2501
rect 2453 -2459 2495 2459
rect 2731 -2459 2773 2459
rect 2453 -2501 2773 -2459
rect -2635 -2740 2429 -2716
rect -2635 -7460 -2611 -2740
rect 2109 -7460 2429 -2740
rect -2635 -7484 2429 -7460
rect -411 -7650 -91 -7484
rect 2109 -7650 2429 -7484
rect 2453 -2641 2773 -2599
rect 2453 -7559 2495 -2641
rect 2731 -7559 2773 -2641
rect 2453 -7601 2773 -7559
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2751 2600 2249 7600
string parameters w 24.0 l 24.0 val 1.17k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
