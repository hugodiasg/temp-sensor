magic
tech sky130A
magscale 1 2
timestamp 1644161670
<< pwell >>
rect -278 -1058 278 1058
<< mvnmos >>
rect -50 -800 50 800
<< mvndiff >>
rect -108 788 -50 800
rect -108 -788 -96 788
rect -62 -788 -50 788
rect -108 -800 -50 -788
rect 50 788 108 800
rect 50 -788 62 788
rect 96 -788 108 788
rect 50 -800 108 -788
<< mvndiffc >>
rect -96 -788 -62 788
rect 62 -788 96 788
<< mvpsubdiff >>
rect -242 1010 242 1022
rect -242 976 -134 1010
rect 134 976 242 1010
rect -242 964 242 976
rect -242 914 -184 964
rect -242 -914 -230 914
rect -196 -914 -184 914
rect 184 914 242 964
rect -242 -964 -184 -914
rect 184 -914 196 914
rect 230 -914 242 914
rect 184 -964 242 -914
rect -242 -976 242 -964
rect -242 -1010 -134 -976
rect 134 -1010 242 -976
rect -242 -1022 242 -1010
<< mvpsubdiffcont >>
rect -134 976 134 1010
rect -230 -914 -196 914
rect 196 -914 230 914
rect -134 -1010 134 -976
<< poly >>
rect -50 872 50 888
rect -50 838 -34 872
rect 34 838 50 872
rect -50 800 50 838
rect -50 -838 50 -800
rect -50 -872 -34 -838
rect 34 -872 50 -838
rect -50 -888 50 -872
<< polycont >>
rect -34 838 34 872
rect -34 -872 34 -838
<< locali >>
rect -230 914 -196 1010
rect 196 914 230 1010
rect -50 838 -34 872
rect 34 838 50 872
rect -96 788 -62 804
rect -96 -804 -62 -788
rect 62 788 96 804
rect 62 -804 96 -788
rect -50 -872 -34 -838
rect 34 -872 50 -838
rect -230 -976 -196 -914
rect 196 -976 230 -914
rect -230 -1010 -134 -976
rect 134 -1010 230 -976
<< viali >>
rect -196 976 -134 1010
rect -134 976 134 1010
rect 134 976 196 1010
rect -34 838 34 872
rect -96 141 -62 771
rect 62 -315 96 315
rect -34 -872 34 -838
<< metal1 >>
rect -208 1010 208 1016
rect -208 976 -196 1010
rect 196 976 208 1010
rect -208 970 208 976
rect -46 872 46 878
rect -46 838 -34 872
rect 34 838 46 872
rect -46 832 46 838
rect -102 771 -56 783
rect -102 141 -96 771
rect -62 141 -56 771
rect -102 129 -56 141
rect 56 315 102 327
rect 56 -315 62 315
rect 96 -315 102 315
rect 56 -327 102 -315
rect -46 -838 46 -832
rect -46 -872 -34 -838
rect 34 -872 46 -838
rect -46 -878 46 -872
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string FIXED_BBOX -213 -993 213 993
string parameters w 8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
string library sky130
<< end >>
