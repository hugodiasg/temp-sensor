magic
tech sky130A
magscale 1 2
timestamp 1669939930
<< nwell >>
rect -860 7020 -268 8658
rect 4280 6720 4872 8658
rect -860 5680 -268 6718
<< pwell >>
rect -820 4960 -228 5580
rect 3840 5180 4432 6500
<< nmos >>
rect -624 5170 -424 5370
rect 4036 5390 4236 6290
<< pmos >>
rect -664 7239 -464 8439
rect 4476 6939 4676 8439
rect -664 5899 -464 6499
<< ndiff >>
rect -682 5358 -624 5370
rect -682 5182 -670 5358
rect -636 5182 -624 5358
rect -682 5170 -624 5182
rect -424 5358 -366 5370
rect -424 5182 -412 5358
rect -378 5182 -366 5358
rect -424 5170 -366 5182
rect 3978 6278 4036 6290
rect 3978 5402 3990 6278
rect 4024 5402 4036 6278
rect 3978 5390 4036 5402
rect 4236 6278 4294 6290
rect 4236 5402 4248 6278
rect 4282 5402 4294 6278
rect 4236 5390 4294 5402
<< pdiff >>
rect -722 8427 -664 8439
rect -722 7251 -710 8427
rect -676 7251 -664 8427
rect -722 7239 -664 7251
rect -464 8427 -406 8439
rect -464 7251 -452 8427
rect -418 7251 -406 8427
rect -464 7239 -406 7251
rect 4418 8427 4476 8439
rect 4418 6951 4430 8427
rect 4464 6951 4476 8427
rect 4418 6939 4476 6951
rect 4676 8427 4734 8439
rect 4676 6951 4688 8427
rect 4722 6951 4734 8427
rect 4676 6939 4734 6951
rect -722 6487 -664 6499
rect -722 5911 -710 6487
rect -676 5911 -664 6487
rect -722 5899 -664 5911
rect -464 6487 -406 6499
rect -464 5911 -452 6487
rect -418 5911 -406 6487
rect -464 5899 -406 5911
<< ndiffc >>
rect -670 5182 -636 5358
rect -412 5182 -378 5358
rect 3990 5402 4024 6278
rect 4248 5402 4282 6278
<< pdiffc >>
rect -710 7251 -676 8427
rect -452 7251 -418 8427
rect 4430 6951 4464 8427
rect 4688 6951 4722 8427
rect -710 5911 -676 6487
rect -452 5911 -418 6487
<< psubdiff >>
rect 3876 6430 3972 6464
rect 4300 6430 4396 6464
rect 3876 6368 3910 6430
rect -784 5510 -688 5544
rect -360 5510 -264 5544
rect -784 5448 -750 5510
rect -298 5448 -264 5510
rect -784 5030 -750 5092
rect 4362 6368 4396 6430
rect 3876 5250 3910 5312
rect 4362 5250 4396 5312
rect 3876 5216 3972 5250
rect 4300 5216 4396 5250
rect -298 5030 -264 5092
rect -784 4996 -688 5030
rect -360 4996 -264 5030
rect -1624 4400 -1600 4540
rect -1400 4400 -1376 4540
<< nsubdiff >>
rect -824 8588 -728 8622
rect -400 8588 -304 8622
rect -824 8526 -790 8588
rect -338 8526 -304 8588
rect -824 7090 -790 7152
rect -338 7090 -304 7152
rect -824 7056 -728 7090
rect -400 7056 -304 7090
rect 4316 8588 4412 8622
rect 4740 8588 4836 8622
rect 4316 8526 4350 8588
rect 4802 8526 4836 8588
rect 4316 6790 4350 6852
rect 4802 6790 4836 6852
rect 4316 6756 4412 6790
rect 4740 6756 4836 6790
rect -824 6648 -728 6682
rect -400 6648 -304 6682
rect -824 6586 -790 6648
rect -338 6586 -304 6648
rect -824 5750 -790 5812
rect -338 5750 -304 5812
rect -824 5716 -728 5750
rect -400 5716 -304 5750
<< psubdiffcont >>
rect 3972 6430 4300 6464
rect -688 5510 -360 5544
rect -784 5092 -750 5448
rect -298 5092 -264 5448
rect 3876 5312 3910 6368
rect 4362 5312 4396 6368
rect 3972 5216 4300 5250
rect -688 4996 -360 5030
rect -1600 4400 -1400 4540
<< nsubdiffcont >>
rect -728 8588 -400 8622
rect -824 7152 -790 8526
rect -338 7152 -304 8526
rect -728 7056 -400 7090
rect 4412 8588 4740 8622
rect 4316 6852 4350 8526
rect 4802 6852 4836 8526
rect 4412 6756 4740 6790
rect -728 6648 -400 6682
rect -824 5812 -790 6586
rect -338 5812 -304 6586
rect -728 5716 -400 5750
<< poly >>
rect -664 8520 -464 8536
rect -664 8486 -648 8520
rect -480 8486 -464 8520
rect -664 8439 -464 8486
rect -664 7192 -464 7239
rect -664 7158 -648 7192
rect -480 7158 -464 7192
rect -664 7142 -464 7158
rect 4476 8520 4676 8536
rect 4476 8486 4492 8520
rect 4660 8486 4676 8520
rect 4476 8439 4676 8486
rect 4476 6892 4676 6939
rect 4476 6858 4492 6892
rect 4660 6858 4676 6892
rect 4476 6842 4676 6858
rect -664 6580 -464 6596
rect -664 6546 -648 6580
rect -480 6546 -464 6580
rect -664 6499 -464 6546
rect -664 5852 -464 5899
rect -664 5818 -648 5852
rect -480 5818 -464 5852
rect -664 5802 -464 5818
rect -624 5442 -424 5458
rect -624 5408 -608 5442
rect -440 5408 -424 5442
rect -624 5370 -424 5408
rect -624 5132 -424 5170
rect -624 5098 -608 5132
rect -440 5098 -424 5132
rect -624 5082 -424 5098
rect 4036 6362 4236 6378
rect 4036 6328 4052 6362
rect 4220 6328 4236 6362
rect 4036 6290 4236 6328
rect 4036 5352 4236 5390
rect 4036 5318 4052 5352
rect 4220 5318 4236 5352
rect 4036 5302 4236 5318
<< polycont >>
rect -648 8486 -480 8520
rect -648 7158 -480 7192
rect 4492 8486 4660 8520
rect 4492 6858 4660 6892
rect -648 6546 -480 6580
rect -648 5818 -480 5852
rect -608 5408 -440 5442
rect -608 5098 -440 5132
rect 4052 6328 4220 6362
rect 4052 5318 4220 5352
<< locali >>
rect -824 8588 -728 8622
rect -400 8588 -304 8622
rect -824 8526 -790 8588
rect -338 8526 -304 8588
rect -664 8486 -648 8520
rect -480 8486 -464 8520
rect -710 8427 -676 8443
rect -710 7235 -676 7251
rect -452 8427 -418 8443
rect -452 7235 -418 7251
rect -664 7158 -648 7192
rect -480 7158 -464 7192
rect -824 7090 -790 7152
rect -338 7090 -304 7152
rect -824 7056 -728 7090
rect -400 7056 -304 7090
rect 4316 8588 4412 8622
rect 4740 8588 4836 8622
rect 4316 8526 4350 8588
rect 4802 8526 4836 8588
rect 4476 8486 4492 8520
rect 4660 8486 4676 8520
rect 4430 8427 4464 8443
rect 4430 6935 4464 6951
rect 4688 8427 4722 8443
rect 4688 6935 4722 6951
rect 4476 6858 4492 6892
rect 4660 6858 4676 6892
rect 4316 6790 4350 6852
rect 4802 6790 4836 6852
rect 4316 6756 4412 6790
rect 4740 6756 4836 6790
rect -824 6648 -728 6682
rect -400 6648 -304 6682
rect -824 6586 -790 6648
rect -338 6586 -304 6648
rect -664 6546 -648 6580
rect -480 6546 -464 6580
rect -710 6487 -676 6503
rect -710 5895 -676 5911
rect -452 6487 -418 6503
rect -452 5895 -418 5911
rect -664 5818 -648 5852
rect -480 5818 -464 5852
rect -824 5750 -790 5812
rect -338 5750 -304 5812
rect -824 5716 -728 5750
rect -400 5716 -304 5750
rect 3876 6430 3972 6464
rect 4300 6430 4396 6464
rect 3876 6368 3910 6430
rect -784 5510 -688 5544
rect -360 5510 -264 5544
rect -784 5448 -750 5510
rect -298 5448 -264 5510
rect -624 5408 -608 5442
rect -440 5408 -424 5442
rect -670 5358 -636 5374
rect -670 5166 -636 5182
rect -412 5358 -378 5374
rect -412 5166 -378 5182
rect -624 5098 -608 5132
rect -440 5098 -424 5132
rect -784 5030 -750 5092
rect 4362 6368 4396 6430
rect 4036 6328 4052 6362
rect 4220 6328 4236 6362
rect 3990 6278 4024 6294
rect 3990 5386 4024 5402
rect 4248 6278 4282 6294
rect 4248 5386 4282 5402
rect 4036 5318 4052 5352
rect 4220 5318 4236 5352
rect 3876 5250 3910 5312
rect 4362 5250 4396 5312
rect 3876 5216 3972 5250
rect 4300 5216 4396 5250
rect -298 5030 -264 5092
rect -784 4996 -688 5030
rect -360 4996 -264 5030
<< viali >>
rect -1620 4400 -1600 4540
rect -1600 4400 -1400 4540
rect -1400 4400 -1380 4540
<< metal1 >>
rect 1040 8860 1240 9060
rect 600 8700 1620 8860
rect 200 8600 340 8620
rect 200 8500 220 8600
rect 320 8500 340 8600
rect 200 8480 340 8500
rect 600 8440 760 8700
rect 1060 8600 1200 8620
rect 1060 8500 1080 8600
rect 1180 8500 1200 8600
rect 1060 8480 1200 8500
rect 400 8280 760 8440
rect 1460 8420 1620 8700
rect 2860 8600 3000 8620
rect 2860 8500 2880 8600
rect 2980 8500 3000 8600
rect 2860 8480 3000 8500
rect 3140 8600 3280 8620
rect 3140 8500 3160 8600
rect 3260 8500 3280 8600
rect 3140 8480 3280 8500
rect 3400 8600 3540 8620
rect 3400 8500 3420 8600
rect 3520 8500 3540 8600
rect 3400 8480 3540 8500
rect 3640 8600 3780 8620
rect 3640 8500 3660 8600
rect 3760 8500 3780 8600
rect 3640 8480 3780 8500
rect 1280 8280 3880 8420
rect 3040 7560 3620 7580
rect -1910 7260 340 7460
rect 40 7160 340 7260
rect 640 7260 1040 7460
rect 3040 7360 4240 7560
rect -1910 6540 380 6740
rect 640 6500 840 7260
rect 4040 6800 4240 7360
rect 4040 6600 5640 6800
rect -1740 5820 -1340 5840
rect -1740 5660 -1520 5820
rect -1360 5660 -1340 5820
rect -1740 5640 -1340 5660
rect -20 5560 160 6480
rect 420 6300 1040 6500
rect 1300 6340 3580 6540
rect 1020 5820 1220 5840
rect 1020 5660 1040 5820
rect 1200 5660 1220 5820
rect 1020 5640 1220 5660
rect -20 5420 1240 5560
rect -20 5200 160 5420
rect 420 5200 1020 5380
rect 1300 5360 1700 6340
rect 4040 6280 4240 6600
rect 3040 6080 4240 6280
rect 1300 5220 1520 5360
rect 1660 5220 1700 5360
rect 1300 5200 1700 5220
rect 2690 5550 3390 5730
rect 2690 5240 2870 5550
rect 630 5050 810 5200
rect 2690 5140 3680 5240
rect 90 4860 1350 5050
rect 2690 4860 2870 5140
rect 4040 5000 4240 6080
rect -1910 4670 2870 4860
rect 3380 4980 4240 5000
rect 3380 4820 3400 4980
rect 3620 4820 4240 4980
rect 3380 4800 4240 4820
rect -1910 4660 2860 4670
rect -1640 4540 -1360 4660
rect -1640 4400 -1620 4540
rect -1380 4400 -1360 4540
rect -1640 4380 -1360 4400
<< via1 >>
rect 220 8500 320 8600
rect 1080 8500 1180 8600
rect 2880 8500 2980 8600
rect 3160 8500 3260 8600
rect 3420 8500 3520 8600
rect 3660 8500 3760 8600
rect -1520 5660 -1360 5820
rect 1040 5660 1200 5820
rect 1520 5220 1660 5360
rect 3400 4820 3620 4980
<< metal2 >>
rect 180 8600 3880 8680
rect 180 8500 220 8600
rect 320 8500 1080 8600
rect 1180 8500 2880 8600
rect 2980 8500 3160 8600
rect 3260 8500 3420 8600
rect 3520 8500 3660 8600
rect 3760 8500 3880 8600
rect 180 8480 3880 8500
rect -1910 5820 1220 5840
rect -1910 5660 -1520 5820
rect -1360 5660 1040 5820
rect 1200 5660 1220 5820
rect -1910 5640 1220 5660
rect 1500 5360 1680 5380
rect 1500 5220 1520 5360
rect 1660 5220 1680 5360
rect 1500 5200 1680 5220
rect 3380 4980 3640 5000
rect 3380 4820 3400 4980
rect 3620 4820 3640 4980
rect 3380 4800 3640 4820
<< via2 >>
rect 1520 5220 1660 5360
rect 3400 4820 3620 4980
<< metal3 >>
rect 1500 5360 1700 5380
rect 1500 5220 1520 5360
rect 1660 5220 1700 5360
rect 1500 4340 1700 5220
rect 3380 4980 3640 5000
rect 3380 4820 3400 4980
rect 3620 4820 3640 4980
rect 3380 4800 3640 4820
<< via3 >>
rect 3400 4820 3620 4980
<< metal4 >>
rect 3380 4980 3640 5000
rect 3380 4820 3400 4980
rect 3620 4820 3640 4980
rect 3380 4180 3640 4820
use sky130_fd_pr__cap_mim_m3_1_2NYK3R  XCC
timestamp 1668740706
transform 1 0 2170 0 1 2340
box -2250 -2200 2249 2200
use sky130_fd_pr__pfet_01v8_G8TFUZ  XM1
timestamp 1668740706
transform 1 0 296 0 1 6199
box -296 -519 296 519
use sky130_fd_pr__pfet_01v8_G8PDUZ  XM2
timestamp 1668741396
transform 1 0 1156 0 1 6199
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_SXTBPF  XM4
timestamp 1668741396
transform 1 0 1157 0 1 5291
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_XABGW3  XM7
timestamp 1668741396
transform 1 0 3345 0 1 5840
box -425 -660 425 660
use sky130_fd_pr__pfet_01v8_8ALGB7  XM8
timestamp 1668740706
transform 1 0 3343 0 1 7689
box -683 -969 683 969
use sky130_fd_pr__nfet_01v8_SXTBPF  sky130_fd_pr__nfet_01v8_SXTBPF_0
timestamp 1668741396
transform 1 0 297 0 1 5291
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_G8TPYT  sky130_fd_pr__pfet_01v8_G8TPYT_0
timestamp 1668740706
transform 1 0 1156 0 1 7839
box -296 -819 296 819
use sky130_fd_pr__pfet_01v8_G8TPYT  sky130_fd_pr__pfet_01v8_G8TPYT_1
timestamp 1668740706
transform 1 0 296 0 1 7839
box -296 -819 296 819
<< labels >>
flabel metal1 1040 8860 1240 9060 0 FreeSans 128 0 0 0 vd
port 0 nsew
flabel metal1 -1740 7260 -1540 7460 0 FreeSans 128 0 0 0 ib
port 2 nsew
flabel metal1 -1740 6540 -1540 6740 0 FreeSans 128 0 0 0 in1
port 3 nsew
flabel metal1 -1740 5640 -1540 5840 0 FreeSans 128 0 0 0 in2
port 4 nsew
flabel metal1 -1740 4660 -1540 4860 0 FreeSans 128 0 0 0 vs
port 1 nsew
flabel metal1 5440 6600 5640 6800 0 FreeSans 128 0 0 0 out
port 5 nsew
<< end >>
