magic
tech sky130A
magscale 1 2
timestamp 1700063261
<< metal4 >>
rect -3349 1539 3349 1580
rect -3349 -1539 3093 1539
rect 3329 -1539 3349 1539
rect -3349 -1580 3349 -1539
<< via4 >>
rect 3093 -1539 3329 1539
<< mimcap2 >>
rect -3269 1460 2731 1500
rect -3269 -1460 -3229 1460
rect 2691 -1460 2731 1460
rect -3269 -1500 2731 -1460
<< mimcap2contact >>
rect -3229 -1460 2691 1460
<< metal5 >>
rect 3051 1539 3371 1581
rect -3253 1460 2715 1484
rect -3253 -1460 -3229 1460
rect 2691 -1460 2715 1460
rect -3253 -1484 2715 -1460
rect 3051 -1539 3093 1539
rect 3329 -1539 3371 1539
rect 3051 -1581 3371 -1539
<< properties >>
string FIXED_BBOX -3349 -1580 2811 1580
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30.0 l 15 val 917.1 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
