** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator_tb-tran.sch
**.subckt ask-modulator_tb-tran
Vdd vd GND 3.3
Vin in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 50ns 100ns)
x1 vd out in GND ask-modulator
**** begin user architecture code


*.tran 0.2n 30n
.tran 0.005n 100n
*.tran 0.3n 400n
*.tran 0.05n 1.3n

.control
destroy all
run
let t=100n
let id =-i(vdd)
plot id
plot in
plot out 3.2950864
*S
let vrms_rlc=sqrt(integ((out-vd)^2)/t)
let vrms_nmos=sqrt(integ(out^2)/t)
let irms=sqrt(integ((-i(vdd))^2)/t)
let srms_rlc=vrms_rlc*irms
let srms_nmos=vrms_nmos*irms
let srms=srms_rlc+srms_nmos
plot srms
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sym # of pins=4
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sch
.subckt ask-modulator  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=23.3 L=23.3 MF=3 m=3
x1 vd out l0
**** begin user architecture code

*X0 out.t2 out.t3 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X1 out in.t0 gnd gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p
*+ ps=1.798e+07u w=0u l=0u
*X2 out.t4 out.t5 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X3 out.t0 out.t1 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 out.n0 out 6.736
R1 out.t1 out.n0 5.23
R2 out out.t1 3.322
R3 out.n1 out.t3 0.472
R4 out.t1 out.n1 0.471
R5 out.n0 out.t2 0.164
R6 out.t4 out.t0 0.066
R7 out.t2 out.t4 0.066
R8 out.n1 out.t5 0.023
R9 in in.t0 448.61
C0 out in 0.05fF
C1 in.t0 gnd 0.46fF
C2 out.t0 gnd 13.53fF
C3 out.t4 gnd 13.57fF
C4 out.t2 gnd 13.79fF
C5 out.n0 gnd 44.65fF $ **FLOATING
C6 out.t5 gnd 6.18fF
C7 out.t3 gnd 8.90fF
C8 out.n1 gnd 3.13fF $ **FLOATING
C9 out.t1 gnd 58.04fF
C10 out gnd 165.23fF
C11 in gnd 5.60fF

**** end user architecture code
XM1 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XR1 out vd gnd sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym # of
*+ pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sch
.subckt l0  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.077n m=1
Cs1 p1 net1 10.78f m=1
Cs2 p2 net2 10.54f m=1
Rs1 net1 GND 41.95 m=1
Rs2 net2 GND 5.649 m=1
R1 p2 net3 4.88 m=1
.ends

.GLOBAL GND
.end
