magic
tech sky130A
magscale 1 2
timestamp 1677666515
<< metal1 >>
rect -8380 25240 -6200 25260
rect -8380 24760 -8360 25240
rect -6260 24760 -6200 25240
rect -8380 24720 -6200 24760
rect -8900 5852 -8200 5920
rect -8902 5148 -6248 5852
rect -8900 5100 -8200 5148
rect -7300 3401 -6500 3500
rect -7301 3199 -6399 3401
rect -8900 -4800 -8200 -4600
rect -8900 -5200 -8300 -4800
rect -7960 -5200 -7950 -4800
rect -8900 -5420 -8200 -5200
rect -7300 -5590 -7100 3199
rect -6600 1140 -6560 1720
rect -5940 1140 -5900 1720
rect -6600 1100 -5900 1140
rect 5000 -700 26350 -500
rect -6755 -1055 4555 -745
rect -6755 -3755 -6445 -1055
rect -6810 -5200 -6800 -4800
rect -6400 -5200 -6390 -4800
rect -7300 -5790 -6500 -5590
rect -7425 -6380 -6500 -6180
rect -8900 -9034 -8200 -8720
rect -7425 -9034 -7225 -6380
rect 4245 -6845 4555 -1055
rect 5000 -3100 5200 -700
rect 14955 -965 17505 -835
rect 14955 -1175 15085 -965
rect 6015 -1305 15085 -1175
rect 6015 -2320 6145 -1305
rect 15500 -1600 17050 -1100
rect 5000 -3300 6100 -3100
rect 6000 -4500 6200 -4000
rect 14515 -4045 14645 -4040
rect 14145 -4355 14855 -4045
rect 5990 -4800 6000 -4500
rect 6200 -4800 6210 -4500
rect 7850 -5220 7860 -4840
rect 8180 -4920 8190 -4840
rect 8180 -5220 8200 -4920
rect 8120 -5240 8200 -5220
rect 14545 -5745 14855 -4355
rect 14545 -6055 14860 -5745
rect 14545 -6365 14855 -6055
rect 15360 -6260 15740 -5660
rect 16290 -6020 16300 -5660
rect 16460 -6020 16470 -5660
rect 16700 -5800 17000 -1600
rect 17375 -2045 17505 -965
rect 21790 -2045 21800 -1940
rect 17185 -2340 21800 -2045
rect 22300 -2340 22310 -1940
rect 17185 -2355 21955 -2340
rect 16690 -6200 16700 -5800
rect 17000 -6200 17010 -5800
rect 14545 -6675 14860 -6365
rect 15350 -6540 15360 -6260
rect 15740 -6540 15750 -6260
rect 17185 -6365 17495 -2355
rect 18100 -3700 19100 -3680
rect 18090 -4000 18100 -3700
rect 18400 -3880 19100 -3700
rect 18400 -4000 18410 -3880
rect 17700 -4655 19055 -4345
rect 26150 -4540 26350 -700
rect 27100 -1980 27680 -1700
rect 26600 -2000 27680 -1980
rect 26590 -2400 26600 -2000
rect 27100 -2740 27680 -2000
rect 17180 -6420 17495 -6365
rect 17180 -6440 17500 -6420
rect 17180 -6660 17200 -6440
rect 17460 -6660 17500 -6440
rect 14545 -6845 14855 -6675
rect 17180 -6680 17500 -6660
rect 17705 -6845 18015 -4655
rect 18090 -5100 18100 -4800
rect 18400 -5100 18410 -4800
rect 4245 -7155 18015 -6845
rect 14545 -7160 14855 -7155
rect 16945 -7160 18015 -7155
rect 17340 -7175 18015 -7160
rect 15360 -7460 15760 -7420
rect -6700 -7525 -6500 -7500
rect -8900 -9234 -7225 -9034
rect -8900 -9540 -8200 -9234
rect -8400 -9685 -7880 -9680
rect -6755 -9685 -6445 -7525
rect 15360 -7640 15380 -7460
rect 15740 -7640 15760 -7460
rect 15360 -7780 15760 -7640
rect 14545 -7800 17455 -7780
rect 14545 -8060 17200 -7800
rect 17420 -8060 17455 -7800
rect 14545 -8090 17455 -8060
rect -4260 -8660 -4060 -8654
rect -4260 -9066 -4060 -9060
rect -3570 -9100 -3560 -8720
rect -3300 -9120 -3240 -9100
rect 14545 -9185 14855 -8090
rect -1835 -9495 14855 -9185
rect -1835 -9685 -1525 -9495
rect -8400 -9700 -1525 -9685
rect -8400 -9980 -8380 -9700
rect -7900 -9980 -1525 -9700
rect -8400 -9995 -1525 -9980
rect 800 -9700 1160 -9680
rect -8400 -10020 -7880 -9995
rect 800 -10080 820 -9700
rect 1140 -10080 1160 -9700
rect 800 -10160 1160 -10080
rect 6005 -10795 6315 -9495
rect 4300 -11700 6300 -11500
rect -1680 -14300 -1480 -13700
rect 4300 -14300 4500 -11700
rect 17705 -12345 18015 -7175
rect 5790 -12600 5800 -12400
rect 6300 -12600 6310 -12400
rect 14345 -12490 18015 -12345
rect 14335 -12600 18015 -12490
rect 14345 -12655 18015 -12600
rect 8010 -13700 8020 -13320
rect 8280 -13720 8340 -13700
rect -1680 -14500 4500 -14300
rect 18100 -15099 18400 -5100
rect 18710 -6580 18720 -6200
rect 19040 -6420 19050 -6200
rect 19070 -6420 19350 -6280
rect 19040 -6580 19350 -6420
rect 18980 -6600 19350 -6580
rect 19070 -13360 19350 -6600
rect 19070 -13640 27200 -13360
rect 17800 -15699 18600 -15099
rect 26920 -15139 27200 -13640
rect 26600 -15719 27640 -15139
<< via1 >>
rect -8360 24760 -6260 25240
rect -8300 -5200 -7960 -4800
rect -6560 1140 -5940 1720
rect -6800 -5200 -6400 -4800
rect 6000 -4800 6200 -4500
rect 7860 -5220 8180 -4840
rect 16300 -6020 16460 -5660
rect 21800 -2340 22300 -1940
rect 16700 -6200 17000 -5800
rect 15360 -6540 15740 -6260
rect 18100 -4000 18400 -3700
rect 26600 -2400 27100 -2000
rect 17200 -6660 17460 -6440
rect 18100 -5100 18400 -4800
rect 15380 -7640 15740 -7460
rect 17200 -8060 17420 -7800
rect -4260 -9060 -4060 -8660
rect -3560 -9100 -3240 -8720
rect -8380 -9980 -7900 -9700
rect 820 -10080 1140 -9700
rect 5800 -12600 6300 -12400
rect 8020 -13700 8340 -13320
rect 18720 -6580 19040 -6200
<< metal2 >>
rect -8380 25240 -6200 25260
rect -8380 24760 -8360 25240
rect -6260 24760 -6200 25240
rect -8380 24720 -6200 24760
rect -6560 1720 -5940 1730
rect -6600 1140 -6560 1720
rect -5940 1140 -5900 1720
rect -6600 1100 -5900 1140
rect 21800 -1940 22300 -1930
rect 21800 -2350 22300 -2340
rect 26600 -2000 27100 -1990
rect 26600 -2410 27100 -2400
rect 18100 -3700 18400 -3690
rect 6000 -4500 6200 -4490
rect -8300 -4800 -7960 -4790
rect -6800 -4800 -6400 -4790
rect -7960 -5200 -6800 -4800
rect -8300 -5210 -7560 -5200
rect -6800 -5210 -6400 -5200
rect -7960 -8660 -7560 -5210
rect -7960 -9060 -4260 -8660
rect -4060 -9060 -4054 -8660
rect -3560 -8720 -3240 -8710
rect -3560 -9110 -3240 -9100
rect 6000 -9300 6200 -4800
rect 18100 -4800 18400 -4000
rect 7860 -4840 8180 -4830
rect 18100 -5110 18400 -5100
rect 7860 -5230 8180 -5220
rect 16280 -5660 16480 -5640
rect 16280 -6020 16300 -5660
rect 16460 -6020 16480 -5660
rect 17700 -5700 19150 -5250
rect 16280 -6040 16480 -6020
rect 16700 -5750 19150 -5700
rect 16700 -5800 18200 -5750
rect 17000 -6200 18200 -5800
rect 18720 -6200 19040 -6190
rect 16700 -6210 17000 -6200
rect 15360 -6260 15760 -6240
rect 15740 -6540 15760 -6260
rect 15360 -7460 15760 -6540
rect 15360 -7640 15380 -7460
rect 15740 -7640 15760 -7460
rect 15360 -7660 15760 -7640
rect 17180 -6440 17500 -6420
rect 17180 -6660 17200 -6440
rect 17460 -6660 17500 -6440
rect 18720 -6590 19040 -6580
rect 17180 -6680 17500 -6660
rect 17180 -7800 17460 -6680
rect 17180 -8060 17200 -7800
rect 17420 -8060 17460 -7800
rect 17180 -8080 17460 -8060
rect 5400 -9500 6200 -9300
rect -8400 -9700 -7880 -9680
rect -8400 -9980 -8380 -9700
rect -7900 -9980 -7880 -9700
rect -8400 -10020 -7880 -9980
rect 800 -9700 1160 -9680
rect 800 -10080 820 -9700
rect 1140 -10080 1160 -9700
rect 800 -10160 1160 -10080
rect 5400 -12400 5600 -9500
rect 5800 -12400 6300 -12390
rect 5400 -12600 5800 -12400
rect 5400 -15099 5600 -12600
rect 5800 -12610 6300 -12600
rect 8020 -13320 8340 -13310
rect 8020 -13710 8340 -13700
rect 5200 -15699 5900 -15099
<< via2 >>
rect -8360 24760 -6260 25240
rect -6560 1140 -5940 1720
rect 21800 -2340 22300 -1940
rect 26600 -2400 27100 -2000
rect -3560 -9100 -3240 -8720
rect 7860 -5220 8180 -4840
rect 16300 -6020 16460 -5660
rect 18720 -6580 19040 -6200
rect -8380 -9980 -7900 -9700
rect 820 -10080 1140 -9700
rect 8020 -13700 8340 -13320
<< metal3 >>
rect -8380 25240 -6200 25260
rect -8400 24760 -8360 25240
rect -6260 24760 -6200 25240
rect -8400 24720 -6200 24760
rect -8400 -9695 -7920 24720
rect -6570 1720 -5930 1725
rect -6600 1140 -6560 1720
rect -5940 1140 -5900 1720
rect -6600 1100 -5900 1140
rect -6410 -590 -6030 1100
rect -6410 -970 4910 -590
rect 4530 -5730 4910 -970
rect 21790 -1940 22310 -1935
rect 21790 -2340 21800 -1940
rect 22300 -2340 22310 -1940
rect 21790 -2345 22310 -2340
rect 26590 -2000 27110 -1995
rect 26590 -2400 26600 -2000
rect 27100 -2400 27110 -2000
rect 26590 -2405 27110 -2400
rect 7840 -4840 8220 -4820
rect 7840 -4880 7860 -4840
rect 7820 -5220 7860 -4880
rect 8180 -5220 8220 -4840
rect 7840 -5730 8220 -5220
rect 4530 -6110 8220 -5730
rect 7840 -6190 8220 -6110
rect 16220 -5660 16560 -5650
rect 16220 -6020 16300 -5660
rect 16460 -6020 16560 -5660
rect 16220 -6190 16560 -6020
rect 7840 -6240 16560 -6190
rect 18710 -6200 19050 -6195
rect 18710 -6240 18720 -6200
rect 7840 -6570 18720 -6240
rect -3640 -8680 -3040 -8580
rect -3640 -8720 1660 -8680
rect -3640 -9100 -3560 -8720
rect -3240 -9100 1660 -8720
rect -3640 -9180 1660 -9100
rect -3600 -9200 1660 -9180
rect 1140 -9600 1660 -9200
rect 640 -9620 1660 -9600
rect 7840 -9620 8220 -6570
rect 16220 -6580 18720 -6570
rect 19040 -6580 19050 -6200
rect 18710 -6585 19050 -6580
rect -8400 -9700 -7890 -9695
rect -8400 -9980 -8380 -9700
rect -7900 -9980 -7890 -9700
rect -8400 -9985 -7890 -9980
rect 640 -9700 8220 -9620
rect -8400 -10020 -7920 -9985
rect 640 -10080 820 -9700
rect 1140 -10080 8220 -9700
rect 640 -10140 8220 -10080
rect 7840 -13300 8220 -10140
rect 7840 -13320 8520 -13300
rect 7840 -13700 8020 -13320
rect 8340 -13700 8520 -13320
rect 7840 -13870 8520 -13700
rect 7860 -13880 8520 -13870
<< via3 >>
rect 21800 -2340 22300 -1940
rect 26600 -2400 27100 -2000
<< metal4 >>
rect 21799 -1940 22301 -1939
rect 21799 -2340 21800 -1940
rect 22300 -2340 22301 -1940
rect 21799 -2341 22301 -2340
rect 26599 -2000 27101 -1999
rect 26599 -2400 26600 -2000
rect 27100 -2400 27101 -2000
rect 26599 -2401 27101 -2400
<< via4 >>
rect 21800 -2340 22300 -1940
rect 26600 -2400 27100 -2000
<< metal5 >>
rect 21776 -1940 22324 -1916
rect 21760 -2340 21800 -1940
rect 22300 -2000 22324 -1940
rect 26576 -2000 27124 -1976
rect 22300 -2340 26600 -2000
rect 21776 -2364 26600 -2340
rect 22000 -2400 26600 -2364
rect 27100 -2400 27124 -2000
rect 26576 -2424 27124 -2400
use ask-modulator  ask-modulator_0 ~/projects-sky130/temp-sensor/ask_modulator/mag
timestamp 1677546845
transform 1 0 -13100 0 1 8600
box 6300 -8800 38800 17562
use buffer  buffer_0 ~/projects-sky130/temp-sensor/buffer/mag
timestamp 1669916246
transform 1 0 -7875 0 1 -6430
box 13875 1430 22120 4938
use buffer  buffer_1
timestamp 1669916246
transform 1 0 -7675 0 1 -14830
box 13875 1430 22120 4938
use ota  ota_0 ~/projects-sky130/temp-sensor/ota/mag
timestamp 1669939930
transform 1 0 20710 0 1 -11140
box -1910 140 5640 9060
use sensor  sensor_0 ~/projects-sky130/temp-sensor/sensor/mag
timestamp 1657129226
transform 1 0 -9100 0 1 -15200
box 2500 1200 11592 5340
use sigma-delta  sigma-delta_0 ~/projects-sky130/temp-sensor/sigma-delta_modulator/mag
timestamp 1675537428
transform 1 0 -1890 0 1 -7930
box -4810 -1070 5739 6386
use sky130_fd_pr__res_xhigh_po_0p35_FT5NBF  sky130_fd_pr__res_xhigh_po_0p35_FT5NBF_0
timestamp 1675991947
transform 1 0 16348 0 1 -3655
box -201 -2598 201 2598
use sky130_fd_pr__res_xhigh_po_0p35_FT5NBF  sky130_fd_pr__res_xhigh_po_0p35_FT5NBF_1
timestamp 1675991947
transform 1 0 15548 0 1 -3655
box -201 -2598 201 2598
<< labels >>
flabel metal1 4400 -12200 4400 -12000 0 FreeSans 1600 0 0 0 vts
flabel metal1 17200 -12500 17200 -12500 0 FreeSans 1600 0 0 0 out_buf1
flabel metal1 8000 -600 8100 -600 0 FreeSans 1600 0 0 0 out_ota
flabel metal1 -7200 -2100 -7200 -2100 0 FreeSans 1600 0 0 0 out_sigma
flabel metal1 -8760 5620 -8740 5620 0 FreeSans 16000 0 0 0 out
port 1 nsew
flabel metal1 -8740 -4960 -8740 -4960 0 FreeSans 16000 0 0 0 vpwr
port 2 nsew
flabel metal1 27420 -2180 27420 -2180 0 FreeSans 16000 0 0 0 vd
port 4 nsew
flabel metal2 5520 -15379 5520 -15379 0 FreeSans 16000 0 0 0 ib2
port 7 nsew
flabel metal1 18220 -15339 18220 -15339 0 FreeSans 16000 0 0 0 ib
port 6 nsew
flabel metal1 27140 -15439 27140 -15439 0 FreeSans 16000 0 0 0 gnd
port 5 nsew
flabel metal1 -8800 -9140 -8680 -9000 0 FreeSans 16000 0 0 0 clk
port 10 nsew
<< end >>
