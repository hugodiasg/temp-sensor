magic
tech sky130A
magscale 1 2
timestamp 1669561651
<< nwell >>
rect -3920 2460 -3610 2720
<< psubdiff >>
rect -1664 -830 -1640 -640
rect -1340 -830 -1316 -640
<< nsubdiff >>
rect -3880 2607 -3853 2641
rect -3695 2607 -3668 2641
<< psubdiffcont >>
rect -1640 -830 -1340 -640
<< nsubdiffcont >>
rect -3853 2607 -3695 2641
<< locali >>
rect -3880 2607 -3853 2641
rect -3695 2607 -3668 2641
rect -1656 -830 -1640 -640
rect -1340 -830 -1324 -640
<< viali >>
rect -3845 2607 -3703 2641
rect -3890 2160 -3840 2200
rect -2110 2160 -2070 2200
rect -1810 2150 -1750 2220
rect -3560 2090 -3510 2130
rect -1640 -830 -1340 -640
<< metal1 >>
rect -3590 5800 -3370 6230
rect -3250 5800 -3030 6230
rect -2930 5790 -2710 6220
rect -2050 5780 -1830 6210
rect -1710 5800 -1490 6230
rect -1400 5790 -1180 6220
rect -4610 4480 -3540 4590
rect -4810 4280 -3540 4480
rect -4610 4160 -3540 4280
rect -3420 4160 -3200 4590
rect -3070 4170 -2850 4600
rect -2760 4530 -2010 4570
rect -2760 4180 -2740 4530
rect -2030 4180 -2010 4530
rect -2760 4160 -2010 4180
rect -1890 4160 -1670 4590
rect -1550 4170 -1330 4600
rect -1230 4140 -920 4580
rect -3015 3905 -1395 4055
rect -4810 3005 -4610 3070
rect -4810 2870 -4485 3005
rect -4610 2540 -4485 2870
rect -3890 2641 -3640 2660
rect -3890 2607 -3845 2641
rect -3703 2607 -3640 2641
rect -3890 2540 -3640 2607
rect -4610 2450 -3640 2540
rect -1545 2575 -1395 3905
rect -1000 3960 -920 4140
rect -1000 3890 -990 3960
rect -920 3890 -910 3960
rect -1545 2570 -415 2575
rect -1545 2430 -590 2570
rect -410 2430 -400 2570
rect -4810 2240 -4610 2340
rect -4810 2230 -4200 2240
rect -1816 2230 -1744 2232
rect -4810 2150 -4300 2230
rect -4210 2150 -4200 2230
rect -1820 2220 -1630 2230
rect -4810 2140 -4200 2150
rect -4030 2200 -3780 2210
rect -4030 2160 -3890 2200
rect -3840 2160 -3780 2200
rect -4030 2140 -3780 2160
rect -2140 2150 -2130 2210
rect -2060 2150 -2050 2210
rect -1820 2150 -1810 2220
rect -1640 2150 -1630 2220
rect -2130 2140 -2060 2150
rect -1820 2140 -1630 2150
rect -4810 1685 -4610 1750
rect -4030 1685 -3960 2140
rect -3590 2060 -3580 2140
rect -3490 2060 -3480 2140
rect -2390 2136 -2320 2140
rect -1816 2138 -1744 2140
rect -2390 2084 -2381 2136
rect -2329 2084 -2320 2136
rect -2390 2070 -2320 2084
rect -4810 1615 -3960 1685
rect -1890 1875 -1740 1950
rect -1545 1875 -1410 2430
rect -600 2425 -415 2430
rect -1890 1725 -1410 1875
rect -1230 1860 -1160 1920
rect -4810 1550 -4610 1615
rect -3530 1400 -1930 1410
rect -3530 1240 -2050 1400
rect -1940 1240 -1930 1400
rect -3530 1230 -1930 1240
rect -4810 400 -4610 410
rect -3530 400 -3350 1230
rect -4810 220 -3350 400
rect -4810 210 -4610 220
rect -1890 -120 -1740 1725
rect -1160 1570 -1070 1610
rect -1160 1430 -1060 1570
rect -960 1430 -950 1570
rect -1160 1420 -1070 1430
rect -1400 1400 -1230 1410
rect -1400 1240 -1390 1400
rect -1280 1240 -1230 1400
rect -1400 1230 -1230 1240
rect -1230 940 -1150 1180
rect -400 980 -290 990
rect -400 940 -390 980
rect -1230 860 -390 940
rect -1230 -60 -1150 860
rect -400 820 -390 860
rect -300 820 -290 980
rect -400 810 -290 820
rect -1890 -280 -1220 -120
rect -1170 -130 -940 -120
rect -1170 -270 -1050 -130
rect -950 -270 -940 -130
rect -1170 -280 -940 -270
rect -2400 -380 -2290 -370
rect -2400 -480 -2390 -380
rect -2300 -480 -2290 -380
rect -2400 -870 -2290 -480
rect -1640 -634 -1480 -280
rect -1220 -380 -1150 -320
rect -1652 -640 -1328 -634
rect -1680 -830 -1640 -640
rect -1340 -830 -1310 -640
rect -1652 -836 -1328 -830
rect -1640 -870 -1480 -836
rect -2450 -1070 -2250 -870
rect -1650 -1070 -1450 -870
<< via1 >>
rect -2740 4180 -2030 4530
rect -990 3890 -920 3960
rect -590 2430 -410 2570
rect -4300 2150 -4210 2230
rect -2130 2200 -2060 2210
rect -2130 2160 -2110 2200
rect -2110 2160 -2070 2200
rect -2070 2160 -2060 2200
rect -2130 2150 -2060 2160
rect -1750 2150 -1640 2220
rect -3580 2130 -3490 2140
rect -3580 2090 -3560 2130
rect -3560 2090 -3510 2130
rect -3510 2090 -3490 2130
rect -3580 2060 -3490 2090
rect -2381 2084 -2329 2136
rect -2050 1240 -1940 1400
rect -1060 1430 -960 1570
rect -1390 1240 -1280 1400
rect -390 820 -300 980
rect -1050 -270 -950 -130
rect -2390 -480 -2300 -380
<< metal2 >>
rect -2760 4530 -2010 4570
rect -2760 4180 -2740 4530
rect -2030 4180 -2010 4530
rect -2760 4160 -2010 4180
rect -2140 3960 -915 3975
rect -2140 3890 -990 3960
rect -920 3890 -915 3960
rect -2140 3885 -915 3890
rect -4310 2230 -4200 2240
rect -4310 2150 -4300 2230
rect -4210 2150 -4200 2230
rect -2140 2210 -2050 3885
rect -990 3880 -920 3885
rect -600 2570 -400 2580
rect -600 2430 -590 2570
rect -410 2430 -400 2570
rect -600 2420 -400 2430
rect -2140 2150 -2130 2210
rect -2060 2150 -2050 2210
rect -4310 2140 -4200 2150
rect -3580 2140 -3490 2150
rect -2140 2140 -2050 2150
rect -1760 2220 -1630 2230
rect -1760 2150 -1750 2220
rect -1640 2150 -1630 2220
rect -1760 2140 -1630 2150
rect -2390 2136 -2320 2140
rect -2390 2084 -2381 2136
rect -2329 2084 -2320 2136
rect -2390 2070 -2320 2084
rect -3580 1685 -3490 2060
rect -3360 1690 -3240 1700
rect -3360 1685 -3350 1690
rect -3580 1595 -3350 1685
rect -3360 1590 -3350 1595
rect -3250 1590 -3240 1690
rect -3360 1580 -3240 1590
rect -2380 -370 -2330 2070
rect -1070 1570 -940 1610
rect -1070 1430 -1060 1570
rect -960 1430 -940 1570
rect -2060 1400 -1270 1410
rect -2060 1240 -2050 1400
rect -1940 1240 -1390 1400
rect -1280 1240 -1270 1400
rect -2060 1230 -1270 1240
rect -1070 740 -940 1430
rect -400 980 -290 990
rect -400 820 -390 980
rect -300 820 -290 980
rect -400 810 -290 820
rect -1060 730 -940 740
rect -1060 650 -1050 730
rect -950 650 -940 730
rect -1060 -130 -940 650
rect -1060 -270 -1050 -130
rect -950 -270 -940 -130
rect -1060 -280 -940 -270
rect -2400 -380 -2290 -370
rect -2400 -480 -2390 -380
rect -2300 -480 -2290 -380
rect -2400 -490 -2290 -480
<< via2 >>
rect -2740 4180 -2030 4530
rect -4300 2150 -4210 2230
rect -590 2430 -410 2570
rect -1750 2150 -1640 2220
rect -3350 1590 -3250 1690
rect -390 820 -300 980
rect -1050 650 -950 730
<< metal3 >>
rect -2760 4530 -2010 4570
rect -2760 4180 -2740 4530
rect -2030 4180 -2010 4530
rect -2760 4160 -2010 4180
rect -600 2570 490 2590
rect -600 2430 -590 2570
rect -410 2430 490 2570
rect -600 2410 490 2430
rect -4310 2230 -1630 2240
rect -4310 2150 -4300 2230
rect -4210 2220 -1630 2230
rect -4210 2150 -1750 2220
rect -1640 2150 -1630 2220
rect -4310 2140 -1630 2150
rect -3360 1690 -3150 1700
rect -3360 1590 -3350 1690
rect -3250 1590 -1530 1690
rect -3360 1580 -3150 1590
rect -1630 740 -1530 1590
rect -400 980 -290 990
rect -400 820 -390 980
rect -300 820 -290 980
rect -400 810 -290 820
rect -1630 730 -940 740
rect -1630 650 -1050 730
rect -950 650 -940 730
rect -1630 640 -940 650
<< via3 >>
rect -2740 4180 -2030 4530
rect -390 820 -300 980
<< metal4 >>
rect -2760 4530 -2010 4570
rect -2760 4180 -2740 4530
rect -2030 4330 -2010 4530
rect -2030 4180 -120 4330
rect -2760 4160 -120 4180
rect -2490 4150 -120 4160
rect -300 990 -120 4150
rect -400 980 340 990
rect -400 820 -390 980
rect -300 820 340 980
rect -400 810 340 820
use sky130_fd_pr__cap_mim_m3_1_A4KLY5  XC1
timestamp 1669420244
transform 1 0 2870 0 1 3420
box -2870 -2820 2869 2820
use sky130_fd_pr__nfet_01v8_X78HBF  XN1
timestamp 1669420244
transform 1 0 -1189 0 1 -190
box -211 -310 211 310
use sky130_fd_pr__res_xhigh_po_0p35_EK42PW  XR2
timestamp 1669420244
transform 1 0 -1614 0 1 5188
box -616 -1198 616 1198
use sky130_fd_pr__pfet_01v8_EFDHR4  sky130_fd_pr__pfet_01v8_EFDHR4_0
timestamp 1669420244
transform 1 0 -1189 0 1 1519
box -211 -519 211 519
use sky130_fd_pr__res_xhigh_po_0p35_ARMGAU  sky130_fd_pr__res_xhigh_po_0p35_ARMGAU_0
timestamp 1669420244
transform 1 0 -3144 0 1 5188
box -616 -1198 616 1198
use sky130_fd_sc_hd__dfrbp_1  x1 ~/sky130_workspace-centos7/open_pdks/sky130/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 -3862 0 1 1948
box -38 -48 2154 592
<< labels >>
flabel metal1 -4810 4280 -4610 4480 0 FreeSans 1600 0 0 0 in
port 1 nsew
flabel metal1 -1650 -1070 -1450 -870 0 FreeSans 1600 0 0 0 gnd
port 6 nsew
flabel metal1 -2450 -1070 -2250 -870 0 FreeSans 1600 0 0 0 reset_b_dff
port 5 nsew
flabel metal1 -4810 1550 -4610 1750 0 FreeSans 1600 0 0 0 clk
port 4 nsew
flabel metal1 -4810 2140 -4610 2340 0 FreeSans 1600 0 0 0 out
port 3 nsew
flabel metal1 -770 890 -720 920 0 FreeSans 800 0 0 0 in_comp
flabel metal3 -1490 670 -1440 700 0 FreeSans 800 0 0 0 out_comp
flabel metal2 -2110 3410 -2080 3470 0 FreeSans 800 0 0 0 Q
flabel metal1 -4810 210 -4610 410 0 FreeSans 1600 0 0 0 vd
port 7 nsew
flabel metal1 -4810 2870 -4610 3070 0 FreeSans 1600 0 0 0 vpwr
port 2 nsew
<< end >>
