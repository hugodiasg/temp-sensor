** sch_path: /foss/designs/temp-sensor/buffer/xschem/buffer-sensor-tb-temp.sch
**.subckt buffer-sensor-tb-temp
VDD vd GND 1.8
Bvts v_lin GND v=-0.00164*temper+1.42962
ibias1 vd ib2 1u
X2 vd vts out ib2 GND buffer-pex
x1 vd vts vtd GND sensor-pex
**** begin user architecture code


.control
destroy all
save all
set color0=white
set color1=black
dc temp -100 300 1
run

plot out-vts
plot out vts
.endc


 .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/temp-sensor/buffer/xschem/buffer-pex.sym # of pins=5
** sym_path: /foss/designs/temp-sensor/buffer/xschem/buffer-pex.sym
** sch_path: /foss/designs/temp-sensor/buffer/xschem/buffer-pex.sch
.subckt buffer-pex vd in out ib gnd
*.iopin vd
*.iopin ib
*.iopin out
*.iopin in
*.iopin gnd
**** begin user architecture code


* NGSPICE file created from buffer.ext - technology: sky130A

*.subckt buffer vd ib out in gnd
X0 vd.t23 a d vd.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 vd.t42 b.t10 out.t9 vd.t41 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2 vd.t21 a d vd.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 out.t8 b.t11 vd.t40 vd.t39 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4 vd.t38 b.t12 out.t7 vd.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 out.t6 b.t13 vd.t1 vd.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X6 c.t9 in.t0 b.t2 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X7 c.t8 in.t1 b.t6 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X8 b.t8 in.t2 c.t7 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X9 b.t5 in.t3 c.t6 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X10 vd.t19 a d vd.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X11 c.t20 out.t20 a gnd.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X12 c.t19 out.t21 a gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X13 out.t10 d gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a a vd.t17 vd.t16 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X15 gnd.t67 d d gnd.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X16 gnd.t65 d d gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X17 d a vd.t15 vd.t14 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X18 vd.t30 vd.t28 vd.t30 vd.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X19 vd.t48 b.t14 out.t5 vd.t47 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X20 d a vd.t13 vd.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 vd.t11 a d vd.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X22 b.t0 in.t4 c.t5 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X23 d d gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X24 d d gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X25 d a vd.t9 vd.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X26 a out.t22 c.t18 gnd.t24 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X27 a out.t23 c.t17 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X28 c.t16 out.t24 a gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X29 a out.t25 c.t15 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X30 a a a gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=2.32 ps=20.6 w=1 l=1
X31 out.t11 d gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X32 gnd.t55 d out.t12 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X33 out.t13 d gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X34 gnd.t51 d out.t14 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X35 gnd.t49 d out.t15 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X36 gnd.t47 d d gnd.t46 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X37 vd.t36 b.t15 out.t4 vd.t35 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X38 c.t4 in.t5 b.t7 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X39 c.t3 in.t6 b.t9 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X40 out.t26 d sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X41 b.t4 in.t7 c.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X42 d d gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X43 vd.t27 vd.t24 vd.t26 vd.t25 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X44 vd.t7 a d vd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X45 c.t14 out.t27 a gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X46 out.t16 d gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X47 gnd.t41 d d gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X48 d d d gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=2.03 ps=18.1 w=1 l=1
X49 d a vd.t5 vd.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X50 vd.t46 b.t16 out.t3 vd.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 out.t2 b.t17 vd.t44 vd.t43 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X52 d a vd.t3 vd.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X53 out.t1 b.t18 vd.t34 vd.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X54 vd.t50 b.t19 out.t0 vd.t49 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X55 b b.t3 vd.t32 vd.t31 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X56 c.t1 in.t8 b.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X57 gnd.t13 ib.t3 ib.t4 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X58 c.t10 ib.t5 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X59 b.t1 in.t9 c.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X60 ib.t2 ib.t0 ib.t1 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X61 d d gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X62 d d gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X63 a a a gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X64 a out.t28 c.t13 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X65 c.t12 out.t29 a gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X66 a out.t30 c.t11 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X67 gnd.t34 d out.t17 gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X68 out.t18 d gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X69 gnd.t30 d out.t19 gnd.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X70 gnd.t28 d d gnd.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
R0 vd.n28 vd.n25 1304.47
R1 vd.n41 vd.n33 1070.68
R2 vd.t41 vd.t31 537.318
R3 vd.t31 vd.t49 526.24
R4 vd.t16 vd.t18 526.24
R5 vd.t14 vd.t16 512.391
R6 vd.t29 vd.t47 357.289
R7 vd.t47 vd.t0 357.289
R8 vd.t0 vd.t37 357.289
R9 vd.t49 vd.t39 357.289
R10 vd.t33 vd.t41 357.289
R11 vd.t45 vd.t33 357.289
R12 vd.t43 vd.t45 357.289
R13 vd.t6 vd.t12 357.289
R14 vd.t12 vd.t10 357.289
R15 vd.t10 vd.t8 357.289
R16 vd.t20 vd.t14 357.289
R17 vd.t4 vd.t20 357.289
R18 vd.t22 vd.t4 357.289
R19 vd.n24 vd.t29 354.529
R20 vd.n31 vd.t6 282.507
R21 vd.n31 vd.t35 254.811
R22 vd.n40 vd.n37 223.625
R23 vd.n34 vd.t2 204.957
R24 vd.n34 vd.t22 152.333
R25 vd.n26 vd.t43 144.024
R26 vd.n33 vd.n28 127.248
R27 vd.n41 vd.n40 117.835
R28 vd.n38 vd.t25 92.7848
R29 vd.n19 vd.t17 29.2512
R30 vd.n14 vd.t7 29.2303
R31 vd.n9 vd.t42 29.2303
R32 vd.n8 vd.t32 29.2303
R33 vd.n1 vd.t27 28.5795
R34 vd.n2 vd.t48 28.57
R35 vd.n0 vd.t3 28.5655
R36 vd.n0 vd.t26 28.5655
R37 vd.n22 vd.t5 28.5655
R38 vd.n22 vd.t23 28.5655
R39 vd.n20 vd.t15 28.5655
R40 vd.n20 vd.t21 28.5655
R41 vd.n17 vd.t9 28.5655
R42 vd.n17 vd.t19 28.5655
R43 vd.n15 vd.t13 28.5655
R44 vd.n15 vd.t11 28.5655
R45 vd.n12 vd.t44 28.5655
R46 vd.n12 vd.t36 28.5655
R47 vd.n10 vd.t34 28.5655
R48 vd.n10 vd.t46 28.5655
R49 vd.n6 vd.t40 28.5655
R50 vd.n6 vd.t50 28.5655
R51 vd.n4 vd.t1 28.5655
R52 vd.n4 vd.t38 28.5655
R53 vd.n1 vd.t24 19.8115
R54 vd.n3 vd.t28 19.8115
R55 vd.n2 vd.t30 14.2847
R56 vd.n5 vd.n3 1.47391
R57 vd vd.n1 1.0363
R58 vd.n8 vd.n7 1.0005
R59 vd.n19 vd.n18 1.0005
R60 vd.n7 vd.n5 0.813
R61 vd.n11 vd.n9 0.813
R62 vd.n18 vd.n16 0.813
R63 vd.n13 vd.n11 0.78175
R64 vd.n16 vd.n14 0.78175
R65 vd.n23 vd.n21 0.78175
R66 vd.n23 vd.n22 0.665316
R67 vd.n21 vd.n20 0.665316
R68 vd.n18 vd.n17 0.665316
R69 vd.n13 vd.n12 0.665316
R70 vd.n11 vd.n10 0.665316
R71 vd.n7 vd.n6 0.665316
R72 vd.n5 vd.n4 0.665316
R73 vd.n14 vd.n13 0.6255
R74 vd.n16 vd.n15 0.611443
R75 vd.n21 vd.n19 0.59425
R76 vd.n42 vd.n23 0.313
R77 vd.n9 vd.n8 0.21925
R78 vd vd.n42 0.0421667
R79 vd.n40 vd.n39 0.0168558
R80 vd.n39 vd.n38 0.0168558
R81 vd.n37 vd.n36 0.00979742
R82 vd.n25 vd.n24 0.00979742
R83 vd.n41 vd.n35 0.0055
R84 vd.n35 vd.n34 0.0055
R85 vd.n3 vd.n2 0.00500317
R86 vd.n1 vd.n0 0.00454578
R87 vd.n28 vd.n27 0.00186586
R88 vd.n27 vd.n26 0.00186586
R89 vd.n33 vd.n32 0.00173262
R90 vd.n32 vd.n31 0.00173262
R91 vd.n30 vd.n29 0.00111631
R92 vd.n31 vd.n30 0.00111631
R93 vd.n42 vd.n41 0.000511142
R94 b.n0 b.t15 40.2461
R95 b.n2 b.t14 40.2461
R96 b b.t3 39.5317
R97 b.n1 b.t10 39.5292
R98 b.n1 b.t18 39.5292
R99 b.n0 b.t16 39.5292
R100 b.n0 b.t17 39.5292
R101 b.n3 b.t19 39.5292
R102 b.n3 b.t11 39.5292
R103 b.n2 b.t12 39.5292
R104 b.n2 b.t13 39.5292
R105 b.n5 b.t6 17.4005
R106 b.n5 b.t5 17.4005
R107 b.n6 b.t7 17.4005
R108 b.n6 b.t4 17.4005
R109 b.n7 b.t2 17.4005
R110 b.n7 b.t8 17.4005
R111 b.n4 b.t9 17.4005
R112 b.n4 b.t0 17.4005
R113 b.n4 b.n5 3.17253
R114 b.n6 b.n7 2.69321
R115 b.n5 b.n6 2.68836
R116 b.t1 b.n4 2.65092
R117 b.n3 b.n2 2.15117
R118 b.n1 b.n0 2.15117
R119 b b.n1 1.49152
R120 b b.t1 0.968485
R121 b b.n3 0.961845
R122 out.n7 out.t4 30.2161
R123 out.n4 out.t0 29.2293
R124 out.n5 out.t9 28.5655
R125 out.n5 out.t1 28.5655
R126 out.n6 out.t3 28.5655
R127 out.n6 out.t2 28.5655
R128 out.n2 out.t7 28.5655
R129 out.n2 out.t8 28.5655
R130 out.n1 out.t5 28.5655
R131 out.n1 out.t6 28.5655
R132 out.n20 out.t20 26.8319
R133 out.n21 out.t27 25.9449
R134 out.n26 out.t30 25.7428
R135 out.n27 out.t21 25.5407
R136 out.n22 out.t28 25.3386
R137 out.n23 out.t29 25.1365
R138 out.n20 out.t22 24.9306
R139 out.n28 out.t25 24.696
R140 out.n25 out.t24 24.5271
R141 out.n24 out.t23 24.1037
R142 out.n0 out.t15 17.4005
R143 out.n0 out.t10 17.4005
R144 out.n10 out.t19 17.4005
R145 out.n10 out.t18 17.4005
R146 out.n11 out.t14 17.4005
R147 out.n11 out.t13 17.4005
R148 out.n12 out.t17 17.4005
R149 out.n12 out.t16 17.4005
R150 out.n13 out.t12 17.4005
R151 out.n13 out.t11 17.4005
R152 out.n14 out.n13 2.74907
R153 out.n17 out.n9 2.41728
R154 out.n24 out.n23 2.30343
R155 out.n22 out.n21 2.29903
R156 out.n28 out.n27 2.2903
R157 out.n26 out.n25 2.25283
R158 out.n16 out.n15 2.1255
R159 out.n15 out.n14 2.1255
R160 out.n29 out.n19 1.97968
R161 out.n18 out.n17 1.83383
R162 out.n3 out.n1 1.74765
R163 out.n19 out.t26 1.69869
R164 out out.n29 1.60362
R165 out.n29 out.n28 1.24394
R166 out.n8 out.n7 1.04217
R167 out.n4 out.n3 1.0005
R168 out.n9 out.n4 0.938
R169 out.n25 out.n24 0.680308
R170 out.n23 out.n22 0.678839
R171 out.n27 out.n26 0.678839
R172 out.n8 out.n5 0.664316
R173 out.n3 out.n2 0.664316
R174 out.n9 out.n8 0.646333
R175 out.n21 out.n20 0.63023
R176 out.n7 out.n6 0.610444
R177 out.n18 out.n0 0.582399
R178 out.n15 out.n11 0.582399
R179 out.n14 out.n12 0.582399
R180 out.n16 out.n10 0.579923
R181 out.n17 out.n16 0.333833
R182 out.n19 out.n18 0.250559
R183 in.n1 in.t6 27.6073
R184 in.n6 in.t7 27.1628
R185 in.n5 in.t5 26.7019
R186 in.n0 in.t8 26.4053
R187 in.n0 in.t9 26.2229
R188 in.n4 in.t3 25.2012
R189 in.n2 in.t4 25.2012
R190 in.n7 in.t0 24.699
R191 in.n3 in.t1 24.699
R192 in.n8 in.t2 24.1526
R193 in in.n8 2.98635
R194 in.n5 in.n4 2.30564
R195 in.n1 in.n0 2.30482
R196 in.n3 in.n2 2.27981
R197 in.n7 in.n6 2.24388
R198 in.n6 in.n5 0.680761
R199 in.n4 in.n3 0.680308
R200 in.n8 in.n7 0.680308
R201 in.n2 in.n1 0.604164
R202 c c.t10 18.4486
R203 c.n17 c.t7 17.4005
R204 c.n17 c.t20 17.4005
R205 c.n13 c.t2 17.4005
R206 c.n13 c.t14 17.4005
R207 c.n11 c.t13 17.4005
R208 c.n11 c.t4 17.4005
R209 c.n9 c.t6 17.4005
R210 c.n9 c.t12 17.4005
R211 c.n7 c.t17 17.4005
R212 c.n7 c.t8 17.4005
R213 c.n5 c.t5 17.4005
R214 c.n5 c.t16 17.4005
R215 c.n3 c.t11 17.4005
R216 c.n3 c.t3 17.4005
R217 c.n1 c.t0 17.4005
R218 c.n1 c.t19 17.4005
R219 c.n0 c.t15 17.4005
R220 c.n0 c.t1 17.4005
R221 c.n15 c.t18 17.4005
R222 c.n15 c.t9 17.4005
R223 c.n2 c.n0 1.87829
R224 c c.n18 1.52139
R225 c.n18 c.n17 1.51465
R226 c.n4 c.n2 1.08383
R227 c.n6 c.n4 1.08383
R228 c.n10 c.n8 1.08383
R229 c.n12 c.n10 1.08383
R230 c.n14 c.n12 1.08383
R231 c.n8 c.n6 1.04217
R232 c.n16 c.n14 1.04217
R233 c.n6 c.n5 0.776026
R234 c.n14 c.n13 0.766495
R235 c.n4 c.n3 0.766495
R236 c.n12 c.n11 0.766495
R237 c.n10 c.n9 0.766495
R238 c.n8 c.n7 0.766495
R239 c.n2 c.n1 0.766495
R240 c.n16 c.n15 0.766495
R241 c.n18 c.n16 0.333833
R242 gnd.n30 gnd.n29 1273.6
R243 gnd.n26 gnd.n23 1260.8
R244 gnd.n51 gnd.n39 1088.88
R245 gnd.t58 gnd.t48 202.462
R246 gnd.t21 gnd.t60 188.337
R247 gnd.t1 gnd.t64 188.337
R248 gnd.t0 gnd.t35 188.337
R249 gnd.t25 gnd.t29 188.337
R250 gnd.t17 gnd.t31 188.337
R251 gnd.t3 gnd.t40 188.337
R252 gnd.t5 gnd.t62 188.337
R253 gnd.t37 gnd.t6 188.337
R254 gnd.t19 gnd.t42 188.337
R255 gnd.t4 gnd.t27 188.337
R256 gnd.t2 gnd.t44 188.337
R257 gnd.t20 gnd.t54 188.337
R258 gnd.t24 gnd.t56 188.337
R259 gnd.t9 gnd.t66 188.337
R260 gnd.n24 gnd.t50 131.835
R261 gnd.t46 gnd.n34 130.267
R262 gnd.t14 gnd.t9 128.696
R263 gnd.t12 gnd.t7 128.696
R264 gnd.n37 gnd.t52 113.002
R265 gnd.n48 gnd.n47 112.218
R266 gnd.n27 gnd.t58 109.079
R267 gnd.n40 gnd.t16 103.585
R268 gnd.n27 gnd.t39 93.3838
R269 gnd.n39 gnd.n26 88.0946
R270 gnd.n37 gnd.t23 75.3349
R271 gnd.t7 gnd.t14 73.7654
R272 gnd.t26 gnd.t12 73.7654
R273 gnd.n47 gnd.n44 62.7792
R274 gnd.n51 gnd.n50 60.3613
R275 gnd.n34 gnd.t8 58.0708
R276 gnd.n40 gnd.t26 25.112
R277 gnd.n19 gnd.t15 17.4005
R278 gnd.n19 gnd.t13 17.4005
R279 gnd.n17 gnd.t57 17.4005
R280 gnd.n17 gnd.t67 17.4005
R281 gnd.n15 gnd.t45 17.4005
R282 gnd.n15 gnd.t55 17.4005
R283 gnd.n13 gnd.t43 17.4005
R284 gnd.n13 gnd.t28 17.4005
R285 gnd.n11 gnd.t38 17.4005
R286 gnd.n11 gnd.t34 17.4005
R287 gnd.n9 gnd.t53 17.4005
R288 gnd.n9 gnd.t47 17.4005
R289 gnd.n7 gnd.t63 17.4005
R290 gnd.n7 gnd.t51 17.4005
R291 gnd.n5 gnd.t32 17.4005
R292 gnd.n5 gnd.t41 17.4005
R293 gnd.n3 gnd.t36 17.4005
R294 gnd.n3 gnd.t30 17.4005
R295 gnd.n1 gnd.t61 17.4005
R296 gnd.n1 gnd.t65 17.4005
R297 gnd.n0 gnd.t59 17.4005
R298 gnd.n0 gnd.t49 17.4005
R299 gnd.t60 gnd.t11 14.1257
R300 gnd.t64 gnd.t21 14.1257
R301 gnd.t35 gnd.t1 14.1257
R302 gnd.t29 gnd.t0 14.1257
R303 gnd.t31 gnd.t25 14.1257
R304 gnd.t40 gnd.t17 14.1257
R305 gnd.t62 gnd.t3 14.1257
R306 gnd.t50 gnd.t5 14.1257
R307 gnd.t52 gnd.t22 14.1257
R308 gnd.t23 gnd.t46 14.1257
R309 gnd.t8 gnd.t37 14.1257
R310 gnd.t6 gnd.t33 14.1257
R311 gnd.t42 gnd.t18 14.1257
R312 gnd.t27 gnd.t19 14.1257
R313 gnd.t44 gnd.t4 14.1257
R314 gnd.t54 gnd.t2 14.1257
R315 gnd.t56 gnd.t20 14.1257
R316 gnd.t66 gnd.t24 14.1257
R317 gnd.n48 gnd.t10 6.27837
R318 gnd.n2 gnd.n0 1.66573
R319 gnd.n20 gnd.n18 1.3755
R320 gnd.n4 gnd.n2 1.08383
R321 gnd.n8 gnd.n6 1.08383
R322 gnd.n10 gnd.n8 1.08383
R323 gnd.n12 gnd.n10 1.08383
R324 gnd.n16 gnd.n14 1.08383
R325 gnd.n18 gnd.n16 1.08383
R326 gnd.n6 gnd.n4 1.04217
R327 gnd.n14 gnd.n12 1.04217
R328 gnd.n18 gnd.n17 0.582399
R329 gnd.n16 gnd.n15 0.582399
R330 gnd.n14 gnd.n13 0.582399
R331 gnd.n12 gnd.n11 0.582399
R332 gnd.n10 gnd.n9 0.582399
R333 gnd.n8 gnd.n7 0.582399
R334 gnd.n6 gnd.n5 0.582399
R335 gnd.n2 gnd.n1 0.582399
R336 gnd.n4 gnd.n3 0.579923
R337 gnd.n20 gnd.n19 0.57713
R338 gnd.n52 gnd.n20 0.392443
R339 gnd.n50 gnd.n49 0.288252
R340 gnd.n49 gnd.n48 0.288252
R341 gnd.n53 gnd.n52 0.101164
R342 gnd.n53 gnd 0.093
R343 gnd gnd.n53 0.0823584
R344 gnd.n43 gnd.n42 0.0425017
R345 gnd.n44 gnd.n43 0.0425017
R346 gnd.n29 gnd.n28 0.0425017
R347 gnd.n28 gnd.n27 0.0425017
R348 gnd.n46 gnd.n45 0.0425017
R349 gnd.n47 gnd.n46 0.0425017
R350 gnd.n23 gnd.n22 0.0425017
R351 gnd.n22 gnd.n21 0.0425017
R352 gnd.n26 gnd.n25 0.00498892
R353 gnd.n25 gnd.n24 0.00498892
R354 gnd.n39 gnd.n38 0.00466542
R355 gnd.n38 gnd.n37 0.00466542
R356 gnd.n31 gnd.n30 0.00271942
R357 gnd.n34 gnd.n31 0.00271942
R358 gnd.n33 gnd.n32 0.00271942
R359 gnd.n34 gnd.n33 0.00271942
R360 gnd.n36 gnd.n35 0.00258271
R361 gnd.n37 gnd.n36 0.00258271
R362 gnd.n51 gnd.n41 0.00190526
R363 gnd.n41 gnd.n40 0.00190526
R364 gnd.n52 gnd.n51 0.000503131
R365 ib.n1 ib.t5 38.0465
R366 ib.n1 ib.t3 37.3602
R367 ib.n3 ib.t0 18.7313
R368 ib.n3 ib.t2 17.409
R369 ib.n0 ib.t4 17.4005
R370 ib.n0 ib.t1 17.4005
R371 ib ib.n4 1.26488
R372 ib.n2 ib.n1 0.239515
R373 ib.n4 ib.n3 0.0163842
R374 ib.n2 ib.n0 0.00444823
R375 ib.n4 ib.n2 0.00358796
C0 in ib 0.0558f
C1 d ib 0.12f
C2 b ib 0.0167f
C3 ib out 0.0112f
C4 ib a 0.0692f
C5 vd c 0.0419f
C6 in vd 0.145f
C7 vd d 1.97f
C8 in c 1.08f
C9 d c 1.32f
C10 b vd 5.7f
C11 vd a 5.74f
C12 vd out 2.13f
C13 in d 0.207f
C14 b c 1.34f
C15 out c 2.02f
C16 c a 3.88f
C17 b in 2.94f
C18 b d 1.04f
C19 in a 0.643f
C20 in out 2.36f
C21 d a 2.4f
C22 d out 40f
C23 vd ib 4.52e-19
C24 b a 0.126f
C25 b out 2.8f
C26 ib c 0.0951f
C27 out a 3.96f
*.ends



**** end user architecture code
.ends


* expanding   symbol:  /foss/designs/temp-sensor/sensor/xschem/sensor-pex.sym # of pins=4
** sym_path: /foss/designs/temp-sensor/sensor/xschem/sensor-pex.sym
** sch_path: /foss/designs/temp-sensor/sensor/xschem/sensor-pex.sch
.subckt sensor-pex vd vts vtd gnd
*.iopin vd
*.opin vts
*.opin vtd
*.iopin gnd
**** begin user architecture code



* NGSPICE file created from sensor.ext - technology: sky130A

*.subckt sensor vd vts vtd gnd
X0 b.t19 vtd c vd.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X1 gnd b.t8 b gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 vtd b.t21 gnd.t40 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 vtd b.t22 gnd.t39 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 gnd.t68 gnd.t66 gnd.t67 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X5 vts.t24 vtd.t12 vtd.t13 vts.t23 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 gnd.t38 b.t23 vtd gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X7 gnd.t37 b.t24 vtd gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X8 vts.t22 vtd.t16 vtd.t17 vts.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X9 gnd b.t6 b gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X10 gnd b.t4 b gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 c vtd.t24 b.t18 vd.t7 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X12 vtd.t15 vtd.t14 vts.t20 vts.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 gnd b.t27 a gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X14 d vtd.t25 vd.t6 vd.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X15 c vtd.t26 b.t17 vd.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 b b.t0 gnd.t30 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X17 gnd.t65 gnd.t63 gnd.t64 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X18 b b.t12 gnd.t29 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X19 gnd.t62 gnd.t60 gnd.t61 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X20 a a vd.t28 vd.t27 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X21 a b.t30 gnd gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X22 a b.t31 gnd gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X23 vd.t26 a a vd.t25 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X24 vtd b.t32 gnd.t24 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X25 vts.t18 vtd.t20 vtd.t21 vts.t17 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 gnd.t59 gnd.t57 gnd.t58 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X27 vd.t20 vd.t17 vd.t19 vd.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X28 b.t16 vtd.t27 c vd.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 vtd b.t33 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X30 gnd.t21 b.t34 vtd gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X31 gnd.t56 gnd.t54 gnd.t55 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X32 c a d vd.t24 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X33 vtd.t19 vtd.t18 vts.t16 vts.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 gnd.t53 gnd.t51 gnd.t52 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X35 gnd.t50 gnd.t47 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X36 vd.t16 vd.t13 vd.t15 vd.t14 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X37 d a c vd.t23 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X38 b b.t14 gnd.t20 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X39 gnd b.t2 b gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X40 vd.t12 vd.t9 vd.t11 vd.t10 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X41 c a d vd.t22 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X42 vtd.t11 vtd.t10 vts.t14 vts.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X43 gnd b.t37 a gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X44 d a c vd.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X45 gnd b.t38 a gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X46 gnd b.t39 a gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X47 b b.t10 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X48 gnd.t46 gnd.t43 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X49 gnd b.t41 vtd gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X50 a b.t42 gnd gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X51 vts.t7 vts.t4 vts.t6 vts.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X52 vts.t12 vtd.t8 vtd.t9 vts.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X53 vd.t2 vtd.t28 vts.t10 vd.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X54 vtd.t23 vtd.t22 vts.t9 vts.t8 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X55 c c c vd.t0 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=1
X56 vts.t3 vts.t0 vts.t2 vts.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X57 a b.t43 gnd gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
R0 vtd.n0 vtd.t25 64.6855
R1 vtd.n5 vtd.t24 64.3461
R2 vtd.n6 vtd.t26 63.6292
R3 vtd.n5 vtd.t27 63.6292
R4 vtd.n15 vtd.t16 63.6292
R5 vtd.n16 vtd.t10 63.6292
R6 vtd.n18 vtd.t20 63.6292
R7 vtd.n19 vtd.t14 63.6292
R8 vtd.n21 vtd.t8 63.6292
R9 vtd.n22 vtd.t18 63.6292
R10 vtd.n24 vtd.t12 63.6292
R11 vtd.n10 vtd.t22 63.6275
R12 vtd.n11 vtd.t23 14.3646
R13 vtd.n15 vtd.t17 14.3555
R14 vtd.n14 vtd.t21 14.283
R15 vtd.n14 vtd.t11 14.283
R16 vtd.n13 vtd.t9 14.283
R17 vtd.n13 vtd.t15 14.283
R18 vtd.n12 vtd.t13 14.283
R19 vtd.n12 vtd.t19 14.283
R20 vtd.n0 vtd.t28 13.7819
R21 vtd.n9 vtd.n8 4.52354
R22 vtd.n4 vtd.n3 4.5005
R23 vtd.n2 vtd.n1 4.5005
R24 vtd.n2 vtd.n0 3.05785
R25 vtd vtd.n27 1.29247
R26 vtd.n27 vtd.n26 0.981502
R27 vtd.n7 vtd.n6 0.792494
R28 vtd.n6 vtd.n5 0.717388
R29 vtd.n27 vtd.n9 0.41175
R30 vtd.n22 vtd.n21 0.134875
R31 vtd.n19 vtd.n18 0.134875
R32 vtd.n16 vtd.n15 0.134875
R33 vtd.n25 vtd.n24 0.0921667
R34 vtd.n24 vtd.n23 0.0676875
R35 vtd.n23 vtd.n22 0.0676875
R36 vtd.n21 vtd.n20 0.0676875
R37 vtd.n20 vtd.n19 0.0676875
R38 vtd.n18 vtd.n17 0.0676875
R39 vtd.n17 vtd.n16 0.0676875
R40 vtd.n11 vtd.n10 0.0516677
R41 vtd.n9 vtd.n4 0.03425
R42 vtd.n4 vtd.n2 0.0255
R43 vtd.n26 vtd.n25 0.022375
R44 vtd.n26 vtd.n11 0.0219082
R45 vtd.n8 vtd.n7 0.00963498
R46 vtd.n17 vtd.n14 0.00576717
R47 vtd.n20 vtd.n13 0.00576717
R48 vtd.n23 vtd.n12 0.00576717
R49 b.t10 b.t12 74.8549
R50 b.t0 b.t10 74.8549
R51 b.t14 b.t0 74.8549
R52 b.t2 b.t4 74.8549
R53 b.t6 b.t2 74.8549
R54 b.t8 b.t6 74.8549
R55 b.t33 b.t22 74.8549
R56 b.t21 b.t33 74.8549
R57 b.t32 b.t21 74.8549
R58 b.t34 b.t24 74.8549
R59 b.t23 b.t34 74.8549
R60 b.t41 b.t23 74.8549
R61 b.t42 b.t31 74.8549
R62 b.t30 b.t42 74.8549
R63 b.t43 b.t30 74.8549
R64 b.t27 b.t38 74.8549
R65 b.t39 b.t27 74.8549
R66 b.t37 b.t39 74.8549
R67 b.n3 b.t37 38.3763
R68 b.n7 b.t14 37.3622
R69 b.n6 b.t8 37.3602
R70 b.n5 b.t32 37.3602
R71 b.n4 b.t41 37.3602
R72 b.n3 b.t43 37.3602
R73 b.n0 b.t18 14.283
R74 b.n0 b.t16 14.283
R75 b.n1 b.t17 14.283
R76 b.n1 b.t19 14.283
R77 b b.n2 2.56613
R78 b b.n7 1.03722
R79 b.n7 b.n6 1.01707
R80 b.n4 b.n3 1.01657
R81 b.n5 b.n4 1.01657
R82 b.n6 b.n5 1.01657
R83 b.n2 b.n0 0.49917
R84 b.n2 b.n1 0.17267
R85 vd.n45 vd.n37 206.306
R86 vd.n17 vd.n14 168.66
R87 vd.t10 vd.n39 156.245
R88 vd.n5 vd.t7 143.697
R89 vd.n43 vd.t27 143.697
R90 vd.n45 vd.n42 126.871
R91 vd.n2 vd.n1 111.421
R92 vd.n15 vd.t4 86.6752
R93 vd.n7 vd.n4 85.0829
R94 vd.n26 vd.n21 79.0593
R95 vd.n27 vd.t14 71.8492
R96 vd.n5 vd.t18 65.0065
R97 vd.n9 vd.t17 63.6934
R98 vd.n32 vd.t13 63.6821
R99 vd.n49 vd.t9 63.6292
R100 vd.n29 vd.n26 63.2476
R101 vd.n15 vd.t8 60.4447
R102 vd.t4 vd.t1 58.1638
R103 vd.t14 vd.t22 58.1638
R104 vd.n24 vd.t5 42.1974
R105 vd.n35 vd.t21 42.1974
R106 vd.n12 vd.t3 28.5119
R107 vd.n40 vd.t10 21.0989
R108 vd.t5 vd.t24 19.3883
R109 vd.n27 vd.t23 17.1073
R110 vd.n31 vd.t6 14.5056
R111 vd.n8 vd.t2 14.472
R112 vd.n31 vd.t15 14.4415
R113 vd.n50 vd.t12 14.4388
R114 vd.n33 vd.t16 14.4153
R115 vd.n10 vd.t19 14.4127
R116 vd.n48 vd.t11 14.4041
R117 vd.n8 vd.t20 14.3878
R118 vd.n47 vd.t28 14.283
R119 vd.n47 vd.t26 14.283
R120 vd.t18 vd.t0 11.4051
R121 vd.n43 vd.t25 3.42187
R122 vd vd.n50 1.79592
R123 vd.n11 vd.n10 0.868662
R124 vd.n48 vd.n47 0.721906
R125 vd.n49 vd.n48 0.608294
R126 vd.n34 vd.n33 0.576317
R127 vd.n18 vd.n11 0.5755
R128 vd.n30 vd.n18 0.488
R129 vd.n46 vd.n34 0.463
R130 vd.n33 vd.n32 0.344245
R131 vd vd.n46 0.2755
R132 vd.n34 vd.n30 0.238
R133 vd.n9 vd.n8 0.129979
R134 vd.n50 vd.n49 0.100468
R135 vd.n32 vd.n31 0.0321654
R136 vd.n4 vd.n3 0.0307238
R137 vd.n3 vd.n2 0.0302348
R138 vd.n10 vd.n9 0.0267443
R139 vd.n42 vd.n41 0.0175052
R140 vd.n41 vd.n40 0.0175052
R141 vd.n21 vd.n20 0.0150968
R142 vd.n20 vd.n19 0.0150968
R143 vd.n14 vd.n13 0.0122827
R144 vd.n13 vd.n12 0.0122827
R145 vd.n37 vd.n36 0.00973799
R146 vd.n36 vd.n35 0.00973799
R147 vd.n17 vd.n16 0.00391284
R148 vd.n16 vd.n15 0.00391284
R149 vd.n29 vd.n28 0.00391284
R150 vd.n28 vd.n27 0.00391284
R151 vd.n45 vd.n44 0.00391284
R152 vd.n44 vd.n43 0.00391284
R153 vd.n7 vd.n6 0.00391284
R154 vd.n6 vd.n5 0.00391284
R155 vd.n39 vd.n38 0.00347027
R156 vd.n1 vd.n0 0.00347027
R157 vd.n26 vd.n25 0.00275116
R158 vd.n25 vd.n24 0.00275116
R159 vd.n24 vd.n23 0.00162558
R160 vd.n23 vd.n22 0.00162558
R161 vd.n18 vd.n17 0.000532663
R162 vd.n30 vd.n29 0.000532663
R163 vd.n46 vd.n45 0.000532663
R164 vd.n11 vd.n7 0.000532663
R165 gnd.n6 gnd.t8 709.494
R166 gnd.n119 gnd.t10 701.865
R167 gnd.t17 gnd.n27 633.203
R168 gnd.n26 gnd.n25 585
R169 gnd.n111 gnd.n110 585
R170 gnd.n116 gnd.n115 585
R171 gnd.n4 gnd.n3 585
R172 gnd.n76 gnd.t2 472.995
R173 gnd.n4 gnd.n2 398.683
R174 gnd.n116 gnd.n114 381.365
R175 gnd.t44 gnd.n5 366.19
R176 gnd.n34 gnd.t22 270.829
R177 gnd.t48 gnd.n118 270.829
R178 gnd.n76 gnd.t0 251.756
R179 gnd.n28 gnd.t17 167.838
R180 gnd.n78 gnd.n75 163.766
R181 gnd.n121 gnd.n111 156.236
R182 gnd.n37 gnd.n36 153.976
R183 gnd.n35 gnd.n30 150.648
R184 gnd.n37 gnd.n26 148.707
R185 gnd.t10 gnd.n117 137.321
R186 gnd.n8 gnd.n4 65.8829
R187 gnd.n113 gnd.n112 57.226
R188 gnd.n34 gnd.n31 49.5887
R189 gnd.n121 gnd.n116 48.5652
R190 gnd.n103 gnd.t47 37.3602
R191 gnd.n106 gnd.t66 37.3602
R192 gnd.n109 gnd.t54 37.3602
R193 gnd.n13 gnd.t63 37.3602
R194 gnd.n16 gnd.t43 37.3602
R195 gnd.n19 gnd.t60 37.3602
R196 gnd.n119 gnd.t48 22.8874
R197 gnd.n10 gnd.t51 18.6812
R198 gnd.n100 gnd.t57 18.6809
R199 gnd.n50 gnd.t24 17.8538
R200 gnd.n21 gnd.t20 17.7911
R201 gnd.n23 gnd.t29 17.4386
R202 gnd.n22 gnd.t9 17.4307
R203 gnd.n21 gnd.t30 17.4235
R204 gnd.n99 gnd.t59 17.405
R205 gnd.n99 gnd.t58 17.405
R206 gnd.n102 gnd.t50 17.405
R207 gnd.n102 gnd.t49 17.405
R208 gnd.n105 gnd.t68 17.405
R209 gnd.n105 gnd.t67 17.405
R210 gnd.n108 gnd.t56 17.405
R211 gnd.n108 gnd.t55 17.405
R212 gnd.n9 gnd.t53 17.405
R213 gnd.n9 gnd.t52 17.405
R214 gnd.n12 gnd.t65 17.405
R215 gnd.n12 gnd.t64 17.405
R216 gnd.n15 gnd.t46 17.405
R217 gnd.n15 gnd.t45 17.405
R218 gnd.n18 gnd.t62 17.405
R219 gnd.n18 gnd.t61 17.405
R220 gnd.n40 gnd.t38 17.4034
R221 gnd.n44 gnd.t40 17.4034
R222 gnd.n52 gnd.t21 17.4034
R223 gnd.n56 gnd.t23 17.4034
R224 gnd.n64 gnd.t37 17.4034
R225 gnd.n67 gnd.t39 17.4034
R226 gnd.n6 gnd.t44 15.2584
R227 gnd.n8 gnd.n7 9.3005
R228 gnd.n7 gnd.n6 9.3005
R229 gnd.n37 gnd.n29 9.3005
R230 gnd.n29 gnd.n28 9.3005
R231 gnd.n78 gnd.n77 9.3005
R232 gnd.n77 gnd.n76 9.3005
R233 gnd.n121 gnd.n120 9.3005
R234 gnd.n120 gnd.n119 9.3005
R235 gnd.n67 gnd.n66 6.38136
R236 gnd.n56 gnd.n55 5.4504
R237 gnd.n64 gnd.n63 5.3168
R238 gnd.n44 gnd.n43 4.92428
R239 gnd.n52 gnd.n51 4.41733
R240 gnd.n40 gnd.n39 3.98894
R241 gnd.n98 gnd.n97 0.624475
R242 gnd.n62 gnd.n50 0.438
R243 gnd.n73 gnd.n62 0.438
R244 gnd.n74 gnd.n73 0.375501
R245 gnd.n22 gnd.n21 0.3755
R246 gnd.n23 gnd.n22 0.3755
R247 gnd.n24 gnd.n23 0.330858
R248 gnd.n24 gnd.n20 0.290469
R249 gnd.n90 gnd.n87 0.287084
R250 gnd.n74 gnd.n38 0.281539
R251 gnd.n89 gnd.n88 0.278696
R252 gnd.n81 gnd.n80 0.278696
R253 gnd.n79 gnd.n74 0.245825
R254 gnd.n123 gnd.n98 0.244548
R255 gnd.n98 gnd.n79 0.180349
R256 gnd.n38 gnd.n24 0.156539
R257 gnd.n94 gnd.n91 0.143628
R258 gnd.n85 gnd.n82 0.143628
R259 gnd.n86 gnd.n85 0.128841
R260 gnd.n49 gnd.n48 0.128341
R261 gnd.n61 gnd.n60 0.128341
R262 gnd.n72 gnd.n71 0.128341
R263 gnd.n95 gnd.n94 0.1255
R264 gnd.n87 gnd.n86 0.0831431
R265 gnd.n97 gnd.n96 0.08175
R266 gnd.n101 gnd.n100 0.073412
R267 gnd.n11 gnd.n10 0.0734113
R268 gnd.n12 gnd.n11 0.0610469
R269 gnd.n13 gnd.n12 0.0610469
R270 gnd.n15 gnd.n14 0.0610469
R271 gnd.n16 gnd.n15 0.0610469
R272 gnd.n18 gnd.n17 0.0610469
R273 gnd.n19 gnd.n18 0.0610469
R274 gnd.n102 gnd.n101 0.0610469
R275 gnd.n103 gnd.n102 0.0610469
R276 gnd.n105 gnd.n104 0.0610469
R277 gnd.n106 gnd.n105 0.0610469
R278 gnd.n108 gnd.n107 0.0610469
R279 gnd.n109 gnd.n108 0.0610469
R280 gnd.n122 gnd.n109 0.0573558
R281 gnd.n20 gnd.n19 0.0573547
R282 gnd.n72 gnd.n68 0.05725
R283 gnd.n72 gnd.n65 0.05725
R284 gnd.n61 gnd.n57 0.051
R285 gnd.n61 gnd.n53 0.051
R286 gnd.n123 gnd.n122 0.0464211
R287 gnd.n49 gnd.n41 0.04475
R288 gnd.n49 gnd.n45 0.04475
R289 gnd.n14 gnd.n13 0.0426875
R290 gnd.n17 gnd.n16 0.0426875
R291 gnd.n104 gnd.n103 0.0426875
R292 gnd.n107 gnd.n106 0.0426875
R293 gnd gnd.n123 0.0415156
R294 gnd.n10 gnd.n9 0.031274
R295 gnd.n100 gnd.n99 0.0312734
R296 gnd.n68 gnd.n67 0.0144748
R297 gnd.n57 gnd.n56 0.0136712
R298 gnd.n48 gnd.n46 0.013
R299 gnd.n48 gnd.n47 0.013
R300 gnd.n45 gnd.n44 0.0127783
R301 gnd.n60 gnd.n58 0.009875
R302 gnd.n60 gnd.n59 0.009875
R303 gnd.n36 gnd.n35 0.0092427
R304 gnd.n35 gnd.n34 0.0092427
R305 gnd.n93 gnd.n92 0.00902273
R306 gnd.n84 gnd.n83 0.00902273
R307 gnd.n114 gnd.n113 0.00883856
R308 gnd.n2 gnd.n1 0.00883856
R309 gnd.n1 gnd.n0 0.00883856
R310 gnd.n65 gnd.n64 0.00867119
R311 gnd.n53 gnd.n52 0.00831404
R312 gnd.n41 gnd.n40 0.00791722
R313 gnd.n71 gnd.n69 0.00675
R314 gnd.n71 gnd.n70 0.00675
R315 gnd.n96 gnd.n90 0.00635717
R316 gnd.n33 gnd.n32 0.00487141
R317 gnd.n34 gnd.n33 0.00487141
R318 gnd.n94 gnd.n93 0.00476136
R319 gnd.n49 gnd.n42 0.00409445
R320 gnd.n61 gnd.n54 0.00393561
R321 gnd.n86 gnd.n81 0.00353363
R322 gnd.n85 gnd.n84 0.00334091
R323 gnd.n122 gnd.n121 0.00152216
R324 gnd.n20 gnd.n8 0.00152195
R325 gnd.n90 gnd.n89 0.00100166
R326 gnd.n38 gnd.n37 0.000522345
R327 gnd.n79 gnd.n78 0.000522345
R328 gnd.n73 gnd.n72 0.000501021
R329 gnd.n62 gnd.n61 0.000501021
R330 gnd.n50 gnd.n49 0.000501021
R331 gnd.n96 gnd.n95 0.000500579
R332 vts.n22 vts.n17 761.601
R333 vts.n23 vts.n22 641.883
R334 vts.t1 vts.t8 333.303
R335 vts.n16 vts.t5 262.014
R336 vts.n26 vts.t1 237.054
R337 vts.t8 vts.t23 229.925
R338 vts.t11 vts.t15 229.925
R339 vts.t19 vts.t17 229.925
R340 vts.t17 vts.t13 229.925
R341 vts.t13 vts.t21 229.925
R342 vts.n20 vts.t11 130.113
R343 vts.n20 vts.t19 99.8129
R344 vts.n11 vts.t0 63.6292
R345 vts.n4 vts.t4 63.6292
R346 vts.n30 vts.n29 37.8314
R347 vts.n12 vts.t10 16.8006
R348 vts.n5 vts.t6 14.4639
R349 vts.n10 vts.t3 14.4362
R350 vts.n13 vts.t2 14.4313
R351 vts.n4 vts.t7 14.3697
R352 vts.n0 vts.t9 14.283
R353 vts.n0 vts.t24 14.283
R354 vts.n1 vts.t16 14.283
R355 vts.n1 vts.t12 14.283
R356 vts.n2 vts.t20 14.283
R357 vts.n2 vts.t18 14.283
R358 vts.n3 vts.t14 14.283
R359 vts.n3 vts.t22 14.283
R360 vts vts.n32 0.88175
R361 vts.n9 vts.n8 0.6455
R362 vts.n8 vts.n7 0.6455
R363 vts.n7 vts.n6 0.6455
R364 vts.n6 vts.n5 0.450361
R365 vts.n10 vts.n9 0.440551
R366 vts.n31 vts.n30 0.369912
R367 vts.n5 vts.n4 0.0741592
R368 vts.n11 vts.n10 0.0682354
R369 vts.n13 vts.n11 0.0634447
R370 vts.n25 vts.n24 0.0431282
R371 vts.n24 vts.n23 0.0426316
R372 vts.n32 vts.n31 0.0305459
R373 vts.n27 vts.n15 0.0180045
R374 vts.n15 vts.n14 0.0175052
R375 vts.n9 vts.n0 0.0129196
R376 vts.n8 vts.n1 0.0129196
R377 vts.n7 vts.n2 0.0129196
R378 vts.n6 vts.n3 0.0129196
R379 vts.n28 vts.n27 0.0111828
R380 vts.n29 vts.n28 0.0106833
R381 vts.n17 vts.n16 0.00559165
R382 vts.n22 vts.n21 0.00192573
R383 vts.n21 vts.n20 0.00192573
R384 vts.n19 vts.n18 0.00192573
R385 vts.n20 vts.n19 0.00192573
R386 vts.n31 vts.n13 0.00106714
R387 vts.n26 vts.n25 0.00100046
R388 vts.n27 vts.n26 0.00100029
R389 vts.n13 vts.n12 0.000503978
C0 a vts 0.543f
C1 vts b 0.972f
C2 vtd vd 3.41f
C3 a c 0.997f
C4 c b 0.55f
C5 vts d 0.248f
C6 a b 0.821f
C7 c d 0.492f
C8 a d 0.588f
C9 d b 0.0152f
C10 vts vd 0.494f
C11 c vd 0.787f
C12 vts vtd 7.5f
C13 c vtd 1.12f
C14 a vd 2.92f
C15 b vd 0.0693f
C16 a vtd 2.14f
C17 vtd b 4.55f
C18 d vd 0.282f
C19 d vtd 0.3f
C20 vts c 0.166f
*.ends



**** end user architecture code
.ends

.GLOBAL GND
.end
