magic
tech sky130A
timestamp 1645128003
<< metal4 >>
rect 25840 20260 26680 25359
<< metal5 >>
rect 21100 29260 30100 30100
rect 21100 28120 28960 28960
rect 21100 21939 21939 28120
rect 22239 26980 27820 27820
rect 22239 23079 23079 26980
rect 23379 25840 26680 26680
rect 23379 24219 24219 25840
rect 25840 24519 26680 25840
rect 26980 24219 27820 26980
rect 23379 23379 27820 24219
rect 28120 23079 28960 28120
rect 22239 22239 28960 23079
rect 29260 21939 30100 29260
rect 21100 21100 30100 21939
<< end >>
