magic
tech sky130A
magscale 1 2
timestamp 1655684427
<< nwell >>
rect -1199 -1019 1199 1019
<< pmos >>
rect -1003 -800 -803 800
rect -745 -800 -545 800
rect -487 -800 -287 800
rect -229 -800 -29 800
rect 29 -800 229 800
rect 287 -800 487 800
rect 545 -800 745 800
rect 803 -800 1003 800
<< pdiff >>
rect -1061 788 -1003 800
rect -1061 -788 -1049 788
rect -1015 -788 -1003 788
rect -1061 -800 -1003 -788
rect -803 788 -745 800
rect -803 -788 -791 788
rect -757 -788 -745 788
rect -803 -800 -745 -788
rect -545 788 -487 800
rect -545 -788 -533 788
rect -499 -788 -487 788
rect -545 -800 -487 -788
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
rect 487 788 545 800
rect 487 -788 499 788
rect 533 -788 545 788
rect 487 -800 545 -788
rect 745 788 803 800
rect 745 -788 757 788
rect 791 -788 803 788
rect 745 -800 803 -788
rect 1003 788 1061 800
rect 1003 -788 1015 788
rect 1049 -788 1061 788
rect 1003 -800 1061 -788
<< pdiffc >>
rect -1049 -788 -1015 788
rect -791 -788 -757 788
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
rect 757 -788 791 788
rect 1015 -788 1049 788
<< nsubdiff >>
rect -1163 949 -1067 983
rect 1067 949 1163 983
rect -1163 887 -1129 949
rect 1129 887 1163 949
rect -1163 -949 -1129 -887
rect 1129 -949 1163 -887
rect -1163 -983 -1067 -949
rect 1067 -983 1163 -949
<< nsubdiffcont >>
rect -1067 949 1067 983
rect -1163 -887 -1129 887
rect 1129 -887 1163 887
rect -1067 -983 1067 -949
<< poly >>
rect -1003 881 -803 897
rect -1003 847 -987 881
rect -819 847 -803 881
rect -1003 800 -803 847
rect -745 881 -545 897
rect -745 847 -729 881
rect -561 847 -545 881
rect -745 800 -545 847
rect -487 881 -287 897
rect -487 847 -471 881
rect -303 847 -287 881
rect -487 800 -287 847
rect -229 881 -29 897
rect -229 847 -213 881
rect -45 847 -29 881
rect -229 800 -29 847
rect 29 881 229 897
rect 29 847 45 881
rect 213 847 229 881
rect 29 800 229 847
rect 287 881 487 897
rect 287 847 303 881
rect 471 847 487 881
rect 287 800 487 847
rect 545 881 745 897
rect 545 847 561 881
rect 729 847 745 881
rect 545 800 745 847
rect 803 881 1003 897
rect 803 847 819 881
rect 987 847 1003 881
rect 803 800 1003 847
rect -1003 -847 -803 -800
rect -1003 -881 -987 -847
rect -819 -881 -803 -847
rect -1003 -897 -803 -881
rect -745 -847 -545 -800
rect -745 -881 -729 -847
rect -561 -881 -545 -847
rect -745 -897 -545 -881
rect -487 -847 -287 -800
rect -487 -881 -471 -847
rect -303 -881 -287 -847
rect -487 -897 -287 -881
rect -229 -847 -29 -800
rect -229 -881 -213 -847
rect -45 -881 -29 -847
rect -229 -897 -29 -881
rect 29 -847 229 -800
rect 29 -881 45 -847
rect 213 -881 229 -847
rect 29 -897 229 -881
rect 287 -847 487 -800
rect 287 -881 303 -847
rect 471 -881 487 -847
rect 287 -897 487 -881
rect 545 -847 745 -800
rect 545 -881 561 -847
rect 729 -881 745 -847
rect 545 -897 745 -881
rect 803 -847 1003 -800
rect 803 -881 819 -847
rect 987 -881 1003 -847
rect 803 -897 1003 -881
<< polycont >>
rect -987 847 -819 881
rect -729 847 -561 881
rect -471 847 -303 881
rect -213 847 -45 881
rect 45 847 213 881
rect 303 847 471 881
rect 561 847 729 881
rect 819 847 987 881
rect -987 -881 -819 -847
rect -729 -881 -561 -847
rect -471 -881 -303 -847
rect -213 -881 -45 -847
rect 45 -881 213 -847
rect 303 -881 471 -847
rect 561 -881 729 -847
rect 819 -881 987 -847
<< locali >>
rect -1163 949 -1067 983
rect 1067 949 1163 983
rect -1163 887 -1129 949
rect 1129 887 1163 949
rect -1003 847 -987 881
rect -819 847 -803 881
rect -745 847 -729 881
rect -561 847 -545 881
rect -487 847 -471 881
rect -303 847 -287 881
rect -229 847 -213 881
rect -45 847 -29 881
rect 29 847 45 881
rect 213 847 229 881
rect 287 847 303 881
rect 471 847 487 881
rect 545 847 561 881
rect 729 847 745 881
rect 803 847 819 881
rect 987 847 1003 881
rect -1049 788 -1015 804
rect -1049 -804 -1015 -788
rect -791 788 -757 804
rect -791 -804 -757 -788
rect -533 788 -499 804
rect -533 -804 -499 -788
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
rect 499 788 533 804
rect 499 -804 533 -788
rect 757 788 791 804
rect 757 -804 791 -788
rect 1015 788 1049 804
rect 1015 -804 1049 -788
rect -1003 -881 -987 -847
rect -819 -881 -803 -847
rect -745 -881 -729 -847
rect -561 -881 -545 -847
rect -487 -881 -471 -847
rect -303 -881 -287 -847
rect -229 -881 -213 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 213 -881 229 -847
rect 287 -881 303 -847
rect 471 -881 487 -847
rect 545 -881 561 -847
rect 729 -881 745 -847
rect 803 -881 819 -847
rect 987 -881 1003 -847
rect -1163 -949 -1129 -887
rect 1129 -949 1163 -887
rect -1163 -983 -1067 -949
rect 1067 -983 1163 -949
<< viali >>
rect -987 847 -819 881
rect -729 847 -561 881
rect -471 847 -303 881
rect -213 847 -45 881
rect 45 847 213 881
rect 303 847 471 881
rect 561 847 729 881
rect 819 847 987 881
rect -1049 141 -1015 771
rect -791 -315 -757 315
rect -533 141 -499 771
rect -275 -315 -241 315
rect -17 141 17 771
rect 241 -315 275 315
rect 499 141 533 771
rect 757 -315 791 315
rect 1015 141 1049 771
rect -987 -881 -819 -847
rect -729 -881 -561 -847
rect -471 -881 -303 -847
rect -213 -881 -45 -847
rect 45 -881 213 -847
rect 303 -881 471 -847
rect 561 -881 729 -847
rect 819 -881 987 -847
<< metal1 >>
rect -999 881 -807 887
rect -999 847 -987 881
rect -819 847 -807 881
rect -999 841 -807 847
rect -741 881 -549 887
rect -741 847 -729 881
rect -561 847 -549 881
rect -741 841 -549 847
rect -483 881 -291 887
rect -483 847 -471 881
rect -303 847 -291 881
rect -483 841 -291 847
rect -225 881 -33 887
rect -225 847 -213 881
rect -45 847 -33 881
rect -225 841 -33 847
rect 33 881 225 887
rect 33 847 45 881
rect 213 847 225 881
rect 33 841 225 847
rect 291 881 483 887
rect 291 847 303 881
rect 471 847 483 881
rect 291 841 483 847
rect 549 881 741 887
rect 549 847 561 881
rect 729 847 741 881
rect 549 841 741 847
rect 807 881 999 887
rect 807 847 819 881
rect 987 847 999 881
rect 807 841 999 847
rect -1055 771 -1009 783
rect -1055 141 -1049 771
rect -1015 141 -1009 771
rect -539 771 -493 783
rect -1055 129 -1009 141
rect -797 315 -751 327
rect -797 -315 -791 315
rect -757 -315 -751 315
rect -539 141 -533 771
rect -499 141 -493 771
rect -23 771 23 783
rect -539 129 -493 141
rect -281 315 -235 327
rect -797 -327 -751 -315
rect -281 -315 -275 315
rect -241 -315 -235 315
rect -23 141 -17 771
rect 17 141 23 771
rect 493 771 539 783
rect -23 129 23 141
rect 235 315 281 327
rect -281 -327 -235 -315
rect 235 -315 241 315
rect 275 -315 281 315
rect 493 141 499 771
rect 533 141 539 771
rect 1009 771 1055 783
rect 493 129 539 141
rect 751 315 797 327
rect 235 -327 281 -315
rect 751 -315 757 315
rect 791 -315 797 315
rect 1009 141 1015 771
rect 1049 141 1055 771
rect 1009 129 1055 141
rect 751 -327 797 -315
rect -999 -847 -807 -841
rect -999 -881 -987 -847
rect -819 -881 -807 -847
rect -999 -887 -807 -881
rect -741 -847 -549 -841
rect -741 -881 -729 -847
rect -561 -881 -549 -847
rect -741 -887 -549 -881
rect -483 -847 -291 -841
rect -483 -881 -471 -847
rect -303 -881 -291 -847
rect -483 -887 -291 -881
rect -225 -847 -33 -841
rect -225 -881 -213 -847
rect -45 -881 -33 -847
rect -225 -887 -33 -881
rect 33 -847 225 -841
rect 33 -881 45 -847
rect 213 -881 225 -847
rect 33 -887 225 -881
rect 291 -847 483 -841
rect 291 -881 303 -847
rect 471 -881 483 -847
rect 291 -887 483 -881
rect 549 -847 741 -841
rect 549 -881 561 -847
rect 729 -881 741 -847
rect 549 -887 741 -881
rect 807 -847 999 -841
rect 807 -881 819 -847
rect 987 -881 999 -847
rect 807 -887 999 -881
<< properties >>
string FIXED_BBOX -1146 -966 1146 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 1.0 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
