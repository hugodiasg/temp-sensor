magic
tech sky130A
magscale 1 2
timestamp 1645148224
<< mvpsubdiff >>
rect -23398 -19130 -23374 -17659
rect -21874 -19130 -21850 -17659
<< mvpsubdiffcont >>
rect -23374 -19130 -21874 -17659
<< locali >>
rect -23390 -19130 -23374 -17659
rect -21874 -19130 -21858 -17659
<< viali >>
rect -23186 -17806 -22020 -17799
rect -23205 -19005 -21999 -17806
<< metal1 >>
rect -24800 11200 -21400 11400
rect -24800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -24800 9800 -21400 10000
rect 9600 -7200 11400 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11400 -7200
rect 9600 -8400 11400 -8200
rect -24800 -17799 -21800 -17600
rect -24800 -17800 -23186 -17799
rect -22020 -17800 -21800 -17799
rect -24800 -17806 -23200 -17800
rect -22000 -17806 -21800 -17800
rect -24800 -19005 -23205 -17806
rect -21999 -19005 -21800 -17806
rect -24800 -19200 -21800 -19005
<< via1 >>
rect -22600 10000 -21600 11200
rect 9800 -8200 10800 -7200
rect -23200 -17806 -23186 -17800
rect -23186 -17806 -22020 -17800
rect -22020 -17806 -22000 -17800
rect -23200 -19000 -22000 -17806
<< metal2 >>
rect -22800 11200 -21400 11400
rect -22800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -22800 9800 -21400 10000
rect 9600 -7200 11000 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect 9600 -8400 11000 -8200
rect -23400 -17800 -21800 -17600
rect -23400 -19000 -23200 -17800
rect -22000 -19000 -21800 -17800
rect -23400 -19200 -21800 -19000
<< via2 >>
rect -22600 10000 -21600 11200
rect 9800 -8200 10800 -7200
rect -23200 -19000 -22000 -17800
<< metal3 >>
rect -22800 11200 -21400 11400
rect -22800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -22800 9800 -21400 10000
rect 9600 -7200 11000 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect 9600 -8400 11000 -8200
rect -23400 -17800 -21800 -17600
rect -23400 -19000 -23200 -17800
rect -22000 -19000 -21800 -17800
rect -23400 -19200 -21800 -19000
<< via3 >>
rect -22600 10000 -21600 11200
rect 9800 -8200 10800 -7200
rect -23200 -19000 -22000 -17800
<< metal4 >>
rect -22800 11200 -21400 11400
rect -22800 10000 -22600 11200
rect -21600 10000 -21400 11200
rect -22800 9800 -21400 10000
rect -23000 -8200 -21600 -3500
rect -18600 -8200 -17200 -4300
rect -12800 -8200 -11400 -4300
rect 2680 -7000 4360 1998
rect -23000 -9600 -11400 -8200
rect 2600 -7200 4400 -7000
rect 2600 -8200 2800 -7200
rect 4200 -8200 4400 -7200
rect 2600 -8400 4400 -8200
rect 9600 -7200 11000 -7000
rect 9600 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect 9600 -8400 11000 -8200
rect -23000 -17600 -21600 -9600
rect -23425 -17800 -21600 -17600
rect -23425 -19000 -23200 -17800
rect -22000 -19000 -21600 -17800
rect -23425 -19233 -21600 -19000
rect -23000 -28200 -21600 -19233
rect -9000 -28200 -7400 -25200
rect -23000 -28400 -7400 -28200
rect -3400 -28400 -1800 -24800
rect 3400 -28400 5000 -25400
rect 9600 -28400 11200 -25400
rect -23000 -29800 11200 -28400
<< via4 >>
rect -22600 10000 -21600 11200
rect 2800 -8200 4200 -7200
rect 9800 -8200 10800 -7200
<< metal5 >>
rect -22840 11200 11200 11480
rect -22840 10000 -22600 11200
rect -21600 10000 11200 11200
rect -22840 9800 11200 10000
rect -22800 6300 -21400 9800
rect -17600 6500 -16200 9800
rect -13200 6400 -11600 9800
rect -6800 7520 8920 9200
rect -6800 -4842 -5122 7520
rect -4522 5240 6640 6920
rect -4522 -2562 -2842 5240
rect -2242 2960 4360 4640
rect -2242 -282 -562 2960
rect 2680 318 4360 2960
rect 4960 -282 6640 5240
rect -2242 -1962 6640 -282
rect 7240 -2562 8920 7520
rect -4522 -4242 8920 -2562
rect 9520 -4842 11200 9800
rect -6800 -6520 11200 -4842
rect -8800 -7200 11000 -7000
rect -8800 -8200 2800 -7200
rect 4200 -8200 9800 -7200
rect 10800 -8200 11000 -7200
rect -8800 -8400 11000 -8200
rect -8800 -11800 -7600 -8400
rect -2600 -11800 -1400 -8400
rect 3600 -11600 4800 -8400
rect 9800 -11800 11000 -8400
use sky130_fd_pr__cap_mim_m3_2_5MQ5FR  sky130_fd_pr__cap_mim_m3_2_5MQ5FR_0
timestamp 1645148224
transform 1 0 -22271 0 1 700
box -2329 -6900 2351 6900
use sky130_fd_pr__cap_mim_m3_2_5MQ5FR  sky130_fd_pr__cap_mim_m3_2_5MQ5FR_1
timestamp 1645148224
transform 1 0 -17271 0 1 700
box -2329 -6900 2351 6900
use sky130_fd_pr__cap_mim_m3_2_5MQ5FR  sky130_fd_pr__cap_mim_m3_2_5MQ5FR_2
timestamp 1645148224
transform 1 0 -12271 0 1 700
box -2329 -6900 2351 6900
use sky130_fd_pr__cap_mim_m3_2_EJYTBJ  sky130_fd_pr__cap_mim_m3_2_EJYTBJ_0
timestamp 1645148224
transform 1 0 -8157 0 1 -18758
box -2843 -8442 2865 8442
use sky130_fd_pr__cap_mim_m3_2_EJYTBJ  sky130_fd_pr__cap_mim_m3_2_EJYTBJ_1
timestamp 1645148224
transform 1 0 -2157 0 1 -18758
box -2843 -8442 2865 8442
use sky130_fd_pr__cap_mim_m3_2_EJYTBJ  sky130_fd_pr__cap_mim_m3_2_EJYTBJ_2
timestamp 1645148224
transform 1 0 3843 0 1 -18758
box -2843 -8442 2865 8442
use sky130_fd_pr__cap_mim_m3_2_EJYTBJ  sky130_fd_pr__cap_mim_m3_2_EJYTBJ_3
timestamp 1645148224
transform 1 0 9843 0 1 -18758
box -2843 -8442 2865 8442
<< labels >>
flabel metal1 11200 -8000 11400 -7800 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 -24800 10400 -24600 10600 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 -24800 -18400 -24600 -18200 0 FreeSans 256 0 0 0 gnd
port 0 nsew
<< end >>
