magic
tech sky130A
magscale 1 2
timestamp 1645715600
<< metal4 >>
rect -2479 7259 2479 7300
rect -2479 2541 2223 7259
rect 2459 2541 2479 7259
rect -2479 2500 2479 2541
rect -2479 2359 2479 2400
rect -2479 -2359 2223 2359
rect 2459 -2359 2479 2359
rect -2479 -2400 2479 -2359
rect -2479 -2541 2479 -2500
rect -2479 -7259 2223 -2541
rect 2459 -7259 2479 -2541
rect -2479 -7300 2479 -7259
<< via4 >>
rect 2223 2541 2459 7259
rect 2223 -2359 2459 2359
rect 2223 -7259 2459 -2541
<< mimcap2 >>
rect -2379 7160 2221 7200
rect -2379 2640 -1887 7160
rect 1729 2640 2221 7160
rect -2379 2600 2221 2640
rect -2379 2260 2221 2300
rect -2379 -2260 -1887 2260
rect 1729 -2260 2221 2260
rect -2379 -2300 2221 -2260
rect -2379 -2640 2221 -2600
rect -2379 -7160 -1887 -2640
rect 1729 -7160 2221 -2640
rect -2379 -7200 2221 -7160
<< mimcap2contact >>
rect -1887 2640 1729 7160
rect -1887 -2260 1729 2260
rect -1887 -7160 1729 -2640
<< metal5 >>
rect -239 7184 81 7350
rect 2181 7259 2501 7350
rect -1911 7160 1753 7184
rect -1911 2640 -1887 7160
rect 1729 2640 1753 7160
rect -1911 2616 1753 2640
rect -239 2284 81 2616
rect 2181 2541 2223 7259
rect 2459 2541 2501 7259
rect 2181 2359 2501 2541
rect -1911 2260 1753 2284
rect -1911 -2260 -1887 2260
rect 1729 -2260 1753 2260
rect -1911 -2284 1753 -2260
rect -239 -2616 81 -2284
rect 2181 -2359 2223 2359
rect 2459 -2359 2501 2359
rect 2181 -2541 2501 -2359
rect -1911 -2640 1753 -2616
rect -1911 -7160 -1887 -2640
rect 1729 -7160 1753 -2640
rect -1911 -7184 1753 -7160
rect -239 -7350 81 -7184
rect 2181 -7259 2223 -2541
rect 2459 -7259 2501 -2541
rect 2181 -7350 2501 -7259
<< properties >>
string FIXED_BBOX -2479 2500 2321 7300
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23 l 23 val 1.075k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
