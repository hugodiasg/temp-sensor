magic
tech sky130A
magscale 1 2
timestamp 1655684427
<< nwell >>
rect -3483 -1019 3483 1019
<< pmos >>
rect -3287 -800 -1687 800
rect -1629 -800 -29 800
rect 29 -800 1629 800
rect 1687 -800 3287 800
<< pdiff >>
rect -3345 788 -3287 800
rect -3345 -788 -3333 788
rect -3299 -788 -3287 788
rect -3345 -800 -3287 -788
rect -1687 788 -1629 800
rect -1687 -788 -1675 788
rect -1641 -788 -1629 788
rect -1687 -800 -1629 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 1629 788 1687 800
rect 1629 -788 1641 788
rect 1675 -788 1687 788
rect 1629 -800 1687 -788
rect 3287 788 3345 800
rect 3287 -788 3299 788
rect 3333 -788 3345 788
rect 3287 -800 3345 -788
<< pdiffc >>
rect -3333 -788 -3299 788
rect -1675 -788 -1641 788
rect -17 -788 17 788
rect 1641 -788 1675 788
rect 3299 -788 3333 788
<< nsubdiff >>
rect -3447 949 -3351 983
rect 3351 949 3447 983
rect -3447 887 -3413 949
rect 3413 887 3447 949
rect -3447 -949 -3413 -887
rect 3413 -949 3447 -887
rect -3447 -983 -3351 -949
rect 3351 -983 3447 -949
<< nsubdiffcont >>
rect -3351 949 3351 983
rect -3447 -887 -3413 887
rect 3413 -887 3447 887
rect -3351 -983 3351 -949
<< poly >>
rect -3287 881 -1687 897
rect -3287 847 -3271 881
rect -1703 847 -1687 881
rect -3287 800 -1687 847
rect -1629 881 -29 897
rect -1629 847 -1613 881
rect -45 847 -29 881
rect -1629 800 -29 847
rect 29 881 1629 897
rect 29 847 45 881
rect 1613 847 1629 881
rect 29 800 1629 847
rect 1687 881 3287 897
rect 1687 847 1703 881
rect 3271 847 3287 881
rect 1687 800 3287 847
rect -3287 -847 -1687 -800
rect -3287 -881 -3271 -847
rect -1703 -881 -1687 -847
rect -3287 -897 -1687 -881
rect -1629 -847 -29 -800
rect -1629 -881 -1613 -847
rect -45 -881 -29 -847
rect -1629 -897 -29 -881
rect 29 -847 1629 -800
rect 29 -881 45 -847
rect 1613 -881 1629 -847
rect 29 -897 1629 -881
rect 1687 -847 3287 -800
rect 1687 -881 1703 -847
rect 3271 -881 3287 -847
rect 1687 -897 3287 -881
<< polycont >>
rect -3271 847 -1703 881
rect -1613 847 -45 881
rect 45 847 1613 881
rect 1703 847 3271 881
rect -3271 -881 -1703 -847
rect -1613 -881 -45 -847
rect 45 -881 1613 -847
rect 1703 -881 3271 -847
<< locali >>
rect -3447 887 -3413 983
rect 3413 887 3447 983
rect -3287 847 -3271 881
rect -1703 847 -1687 881
rect -1629 847 -1613 881
rect -45 847 -29 881
rect 29 847 45 881
rect 1613 847 1629 881
rect 1687 847 1703 881
rect 3271 847 3287 881
rect -3333 788 -3299 804
rect -3333 -804 -3299 -788
rect -1675 788 -1641 804
rect -1675 -804 -1641 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 1641 788 1675 804
rect 1641 -804 1675 -788
rect 3299 788 3333 804
rect 3299 -804 3333 -788
rect -3287 -881 -3271 -847
rect -1703 -881 -1687 -847
rect -1629 -881 -1613 -847
rect -45 -881 -29 -847
rect 29 -881 45 -847
rect 1613 -881 1629 -847
rect 1687 -881 1703 -847
rect 3271 -881 3287 -847
rect -3447 -949 -3413 -887
rect 3413 -949 3447 -887
rect -3447 -983 -3351 -949
rect 3351 -983 3447 -949
<< viali >>
rect -3413 949 -3351 983
rect -3351 949 3351 983
rect 3351 949 3413 983
rect -3271 847 -1703 881
rect -1613 847 -45 881
rect 45 847 1613 881
rect 1703 847 3271 881
rect -3333 141 -3299 771
rect -1675 -315 -1641 315
rect -17 141 17 771
rect 1641 -315 1675 315
rect 3299 141 3333 771
rect -3271 -881 -1703 -847
rect -1613 -881 -45 -847
rect 45 -881 1613 -847
rect 1703 -881 3271 -847
<< metal1 >>
rect -3425 983 3425 989
rect -3425 949 -3413 983
rect 3413 949 3425 983
rect -3425 943 3425 949
rect -3283 881 -1691 887
rect -3283 847 -3271 881
rect -1703 847 -1691 881
rect -3283 841 -1691 847
rect -1625 881 -33 887
rect -1625 847 -1613 881
rect -45 847 -33 881
rect -1625 841 -33 847
rect 33 881 1625 887
rect 33 847 45 881
rect 1613 847 1625 881
rect 33 841 1625 847
rect 1691 881 3283 887
rect 1691 847 1703 881
rect 3271 847 3283 881
rect 1691 841 3283 847
rect -3339 771 -3293 783
rect -3339 141 -3333 771
rect -3299 141 -3293 771
rect -23 771 23 783
rect -3339 129 -3293 141
rect -1681 315 -1635 327
rect -1681 -315 -1675 315
rect -1641 -315 -1635 315
rect -23 141 -17 771
rect 17 141 23 771
rect 3293 771 3339 783
rect -23 129 23 141
rect 1635 315 1681 327
rect -1681 -327 -1635 -315
rect 1635 -315 1641 315
rect 1675 -315 1681 315
rect 3293 141 3299 771
rect 3333 141 3339 771
rect 3293 129 3339 141
rect 1635 -327 1681 -315
rect -3283 -847 -1691 -841
rect -3283 -881 -3271 -847
rect -1703 -881 -1691 -847
rect -3283 -887 -1691 -881
rect -1625 -847 -33 -841
rect -1625 -881 -1613 -847
rect -45 -881 -33 -847
rect -1625 -887 -33 -881
rect 33 -847 1625 -841
rect 33 -881 45 -847
rect 1613 -881 1625 -847
rect 33 -887 1625 -881
rect 1691 -847 3283 -841
rect 1691 -881 1703 -847
rect 3271 -881 3283 -847
rect 1691 -887 3283 -881
<< properties >>
string FIXED_BBOX -3430 -966 3430 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 8.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
