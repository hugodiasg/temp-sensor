magic
tech sky130A
magscale 1 2
timestamp 1675896495
<< metal4 >>
rect -2669 62839 2669 62880
rect -2669 58121 2413 62839
rect 2649 58121 2669 62839
rect -2669 58080 2669 58121
rect -2669 57799 2669 57840
rect -2669 53081 2413 57799
rect 2649 53081 2669 57799
rect -2669 53040 2669 53081
rect -2669 52759 2669 52800
rect -2669 48041 2413 52759
rect 2649 48041 2669 52759
rect -2669 48000 2669 48041
rect -2669 47719 2669 47760
rect -2669 43001 2413 47719
rect 2649 43001 2669 47719
rect -2669 42960 2669 43001
rect -2669 42679 2669 42720
rect -2669 37961 2413 42679
rect 2649 37961 2669 42679
rect -2669 37920 2669 37961
rect -2669 37639 2669 37680
rect -2669 32921 2413 37639
rect 2649 32921 2669 37639
rect -2669 32880 2669 32921
rect -2669 32599 2669 32640
rect -2669 27881 2413 32599
rect 2649 27881 2669 32599
rect -2669 27840 2669 27881
rect -2669 27559 2669 27600
rect -2669 22841 2413 27559
rect 2649 22841 2669 27559
rect -2669 22800 2669 22841
rect -2669 22519 2669 22560
rect -2669 17801 2413 22519
rect 2649 17801 2669 22519
rect -2669 17760 2669 17801
rect -2669 17479 2669 17520
rect -2669 12761 2413 17479
rect 2649 12761 2669 17479
rect -2669 12720 2669 12761
rect -2669 12439 2669 12480
rect -2669 7721 2413 12439
rect 2649 7721 2669 12439
rect -2669 7680 2669 7721
rect -2669 7399 2669 7440
rect -2669 2681 2413 7399
rect 2649 2681 2669 7399
rect -2669 2640 2669 2681
rect -2669 2359 2669 2400
rect -2669 -2359 2413 2359
rect 2649 -2359 2669 2359
rect -2669 -2400 2669 -2359
rect -2669 -2681 2669 -2640
rect -2669 -7399 2413 -2681
rect 2649 -7399 2669 -2681
rect -2669 -7440 2669 -7399
rect -2669 -7721 2669 -7680
rect -2669 -12439 2413 -7721
rect 2649 -12439 2669 -7721
rect -2669 -12480 2669 -12439
rect -2669 -12761 2669 -12720
rect -2669 -17479 2413 -12761
rect 2649 -17479 2669 -12761
rect -2669 -17520 2669 -17479
rect -2669 -17801 2669 -17760
rect -2669 -22519 2413 -17801
rect 2649 -22519 2669 -17801
rect -2669 -22560 2669 -22519
rect -2669 -22841 2669 -22800
rect -2669 -27559 2413 -22841
rect 2649 -27559 2669 -22841
rect -2669 -27600 2669 -27559
rect -2669 -27881 2669 -27840
rect -2669 -32599 2413 -27881
rect 2649 -32599 2669 -27881
rect -2669 -32640 2669 -32599
rect -2669 -32921 2669 -32880
rect -2669 -37639 2413 -32921
rect 2649 -37639 2669 -32921
rect -2669 -37680 2669 -37639
rect -2669 -37961 2669 -37920
rect -2669 -42679 2413 -37961
rect 2649 -42679 2669 -37961
rect -2669 -42720 2669 -42679
rect -2669 -43001 2669 -42960
rect -2669 -47719 2413 -43001
rect 2649 -47719 2669 -43001
rect -2669 -47760 2669 -47719
rect -2669 -48041 2669 -48000
rect -2669 -52759 2413 -48041
rect 2649 -52759 2669 -48041
rect -2669 -52800 2669 -52759
rect -2669 -53081 2669 -53040
rect -2669 -57799 2413 -53081
rect 2649 -57799 2669 -53081
rect -2669 -57840 2669 -57799
rect -2669 -58121 2669 -58080
rect -2669 -62839 2413 -58121
rect 2649 -62839 2669 -58121
rect -2669 -62880 2669 -62839
<< via4 >>
rect 2413 58121 2649 62839
rect 2413 53081 2649 57799
rect 2413 48041 2649 52759
rect 2413 43001 2649 47719
rect 2413 37961 2649 42679
rect 2413 32921 2649 37639
rect 2413 27881 2649 32599
rect 2413 22841 2649 27559
rect 2413 17801 2649 22519
rect 2413 12761 2649 17479
rect 2413 7721 2649 12439
rect 2413 2681 2649 7399
rect 2413 -2359 2649 2359
rect 2413 -7399 2649 -2681
rect 2413 -12439 2649 -7721
rect 2413 -17479 2649 -12761
rect 2413 -22519 2649 -17801
rect 2413 -27559 2649 -22841
rect 2413 -32599 2649 -27881
rect 2413 -37639 2649 -32921
rect 2413 -42679 2649 -37961
rect 2413 -47719 2649 -43001
rect 2413 -52759 2649 -48041
rect 2413 -57799 2649 -53081
rect 2413 -62839 2649 -58121
<< mimcap2 >>
rect -2589 62760 2051 62800
rect -2589 58200 -2549 62760
rect 2011 58200 2051 62760
rect -2589 58160 2051 58200
rect -2589 57720 2051 57760
rect -2589 53160 -2549 57720
rect 2011 53160 2051 57720
rect -2589 53120 2051 53160
rect -2589 52680 2051 52720
rect -2589 48120 -2549 52680
rect 2011 48120 2051 52680
rect -2589 48080 2051 48120
rect -2589 47640 2051 47680
rect -2589 43080 -2549 47640
rect 2011 43080 2051 47640
rect -2589 43040 2051 43080
rect -2589 42600 2051 42640
rect -2589 38040 -2549 42600
rect 2011 38040 2051 42600
rect -2589 38000 2051 38040
rect -2589 37560 2051 37600
rect -2589 33000 -2549 37560
rect 2011 33000 2051 37560
rect -2589 32960 2051 33000
rect -2589 32520 2051 32560
rect -2589 27960 -2549 32520
rect 2011 27960 2051 32520
rect -2589 27920 2051 27960
rect -2589 27480 2051 27520
rect -2589 22920 -2549 27480
rect 2011 22920 2051 27480
rect -2589 22880 2051 22920
rect -2589 22440 2051 22480
rect -2589 17880 -2549 22440
rect 2011 17880 2051 22440
rect -2589 17840 2051 17880
rect -2589 17400 2051 17440
rect -2589 12840 -2549 17400
rect 2011 12840 2051 17400
rect -2589 12800 2051 12840
rect -2589 12360 2051 12400
rect -2589 7800 -2549 12360
rect 2011 7800 2051 12360
rect -2589 7760 2051 7800
rect -2589 7320 2051 7360
rect -2589 2760 -2549 7320
rect 2011 2760 2051 7320
rect -2589 2720 2051 2760
rect -2589 2280 2051 2320
rect -2589 -2280 -2549 2280
rect 2011 -2280 2051 2280
rect -2589 -2320 2051 -2280
rect -2589 -2760 2051 -2720
rect -2589 -7320 -2549 -2760
rect 2011 -7320 2051 -2760
rect -2589 -7360 2051 -7320
rect -2589 -7800 2051 -7760
rect -2589 -12360 -2549 -7800
rect 2011 -12360 2051 -7800
rect -2589 -12400 2051 -12360
rect -2589 -12840 2051 -12800
rect -2589 -17400 -2549 -12840
rect 2011 -17400 2051 -12840
rect -2589 -17440 2051 -17400
rect -2589 -17880 2051 -17840
rect -2589 -22440 -2549 -17880
rect 2011 -22440 2051 -17880
rect -2589 -22480 2051 -22440
rect -2589 -22920 2051 -22880
rect -2589 -27480 -2549 -22920
rect 2011 -27480 2051 -22920
rect -2589 -27520 2051 -27480
rect -2589 -27960 2051 -27920
rect -2589 -32520 -2549 -27960
rect 2011 -32520 2051 -27960
rect -2589 -32560 2051 -32520
rect -2589 -33000 2051 -32960
rect -2589 -37560 -2549 -33000
rect 2011 -37560 2051 -33000
rect -2589 -37600 2051 -37560
rect -2589 -38040 2051 -38000
rect -2589 -42600 -2549 -38040
rect 2011 -42600 2051 -38040
rect -2589 -42640 2051 -42600
rect -2589 -43080 2051 -43040
rect -2589 -47640 -2549 -43080
rect 2011 -47640 2051 -43080
rect -2589 -47680 2051 -47640
rect -2589 -48120 2051 -48080
rect -2589 -52680 -2549 -48120
rect 2011 -52680 2051 -48120
rect -2589 -52720 2051 -52680
rect -2589 -53160 2051 -53120
rect -2589 -57720 -2549 -53160
rect 2011 -57720 2051 -53160
rect -2589 -57760 2051 -57720
rect -2589 -58200 2051 -58160
rect -2589 -62760 -2549 -58200
rect 2011 -62760 2051 -58200
rect -2589 -62800 2051 -62760
<< mimcap2contact >>
rect -2549 58200 2011 62760
rect -2549 53160 2011 57720
rect -2549 48120 2011 52680
rect -2549 43080 2011 47640
rect -2549 38040 2011 42600
rect -2549 33000 2011 37560
rect -2549 27960 2011 32520
rect -2549 22920 2011 27480
rect -2549 17880 2011 22440
rect -2549 12840 2011 17400
rect -2549 7800 2011 12360
rect -2549 2760 2011 7320
rect -2549 -2280 2011 2280
rect -2549 -7320 2011 -2760
rect -2549 -12360 2011 -7800
rect -2549 -17400 2011 -12840
rect -2549 -22440 2011 -17880
rect -2549 -27480 2011 -22920
rect -2549 -32520 2011 -27960
rect -2549 -37560 2011 -33000
rect -2549 -42600 2011 -38040
rect -2549 -47640 2011 -43080
rect -2549 -52680 2011 -48120
rect -2549 -57720 2011 -53160
rect -2549 -62760 2011 -58200
<< metal5 >>
rect -429 62784 -109 63000
rect 2371 62839 2691 63000
rect -2573 62760 2035 62784
rect -2573 58200 -2549 62760
rect 2011 58200 2035 62760
rect -2573 58176 2035 58200
rect -429 57744 -109 58176
rect 2371 58121 2413 62839
rect 2649 58121 2691 62839
rect 2371 57799 2691 58121
rect -2573 57720 2035 57744
rect -2573 53160 -2549 57720
rect 2011 53160 2035 57720
rect -2573 53136 2035 53160
rect -429 52704 -109 53136
rect 2371 53081 2413 57799
rect 2649 53081 2691 57799
rect 2371 52759 2691 53081
rect -2573 52680 2035 52704
rect -2573 48120 -2549 52680
rect 2011 48120 2035 52680
rect -2573 48096 2035 48120
rect -429 47664 -109 48096
rect 2371 48041 2413 52759
rect 2649 48041 2691 52759
rect 2371 47719 2691 48041
rect -2573 47640 2035 47664
rect -2573 43080 -2549 47640
rect 2011 43080 2035 47640
rect -2573 43056 2035 43080
rect -429 42624 -109 43056
rect 2371 43001 2413 47719
rect 2649 43001 2691 47719
rect 2371 42679 2691 43001
rect -2573 42600 2035 42624
rect -2573 38040 -2549 42600
rect 2011 38040 2035 42600
rect -2573 38016 2035 38040
rect -429 37584 -109 38016
rect 2371 37961 2413 42679
rect 2649 37961 2691 42679
rect 2371 37639 2691 37961
rect -2573 37560 2035 37584
rect -2573 33000 -2549 37560
rect 2011 33000 2035 37560
rect -2573 32976 2035 33000
rect -429 32544 -109 32976
rect 2371 32921 2413 37639
rect 2649 32921 2691 37639
rect 2371 32599 2691 32921
rect -2573 32520 2035 32544
rect -2573 27960 -2549 32520
rect 2011 27960 2035 32520
rect -2573 27936 2035 27960
rect -429 27504 -109 27936
rect 2371 27881 2413 32599
rect 2649 27881 2691 32599
rect 2371 27559 2691 27881
rect -2573 27480 2035 27504
rect -2573 22920 -2549 27480
rect 2011 22920 2035 27480
rect -2573 22896 2035 22920
rect -429 22464 -109 22896
rect 2371 22841 2413 27559
rect 2649 22841 2691 27559
rect 2371 22519 2691 22841
rect -2573 22440 2035 22464
rect -2573 17880 -2549 22440
rect 2011 17880 2035 22440
rect -2573 17856 2035 17880
rect -429 17424 -109 17856
rect 2371 17801 2413 22519
rect 2649 17801 2691 22519
rect 2371 17479 2691 17801
rect -2573 17400 2035 17424
rect -2573 12840 -2549 17400
rect 2011 12840 2035 17400
rect -2573 12816 2035 12840
rect -429 12384 -109 12816
rect 2371 12761 2413 17479
rect 2649 12761 2691 17479
rect 2371 12439 2691 12761
rect -2573 12360 2035 12384
rect -2573 7800 -2549 12360
rect 2011 7800 2035 12360
rect -2573 7776 2035 7800
rect -429 7344 -109 7776
rect 2371 7721 2413 12439
rect 2649 7721 2691 12439
rect 2371 7399 2691 7721
rect -2573 7320 2035 7344
rect -2573 2760 -2549 7320
rect 2011 2760 2035 7320
rect -2573 2736 2035 2760
rect -429 2304 -109 2736
rect 2371 2681 2413 7399
rect 2649 2681 2691 7399
rect 2371 2359 2691 2681
rect -2573 2280 2035 2304
rect -2573 -2280 -2549 2280
rect 2011 -2280 2035 2280
rect -2573 -2304 2035 -2280
rect -429 -2736 -109 -2304
rect 2371 -2359 2413 2359
rect 2649 -2359 2691 2359
rect 2371 -2681 2691 -2359
rect -2573 -2760 2035 -2736
rect -2573 -7320 -2549 -2760
rect 2011 -7320 2035 -2760
rect -2573 -7344 2035 -7320
rect -429 -7776 -109 -7344
rect 2371 -7399 2413 -2681
rect 2649 -7399 2691 -2681
rect 2371 -7721 2691 -7399
rect -2573 -7800 2035 -7776
rect -2573 -12360 -2549 -7800
rect 2011 -12360 2035 -7800
rect -2573 -12384 2035 -12360
rect -429 -12816 -109 -12384
rect 2371 -12439 2413 -7721
rect 2649 -12439 2691 -7721
rect 2371 -12761 2691 -12439
rect -2573 -12840 2035 -12816
rect -2573 -17400 -2549 -12840
rect 2011 -17400 2035 -12840
rect -2573 -17424 2035 -17400
rect -429 -17856 -109 -17424
rect 2371 -17479 2413 -12761
rect 2649 -17479 2691 -12761
rect 2371 -17801 2691 -17479
rect -2573 -17880 2035 -17856
rect -2573 -22440 -2549 -17880
rect 2011 -22440 2035 -17880
rect -2573 -22464 2035 -22440
rect -429 -22896 -109 -22464
rect 2371 -22519 2413 -17801
rect 2649 -22519 2691 -17801
rect 2371 -22841 2691 -22519
rect -2573 -22920 2035 -22896
rect -2573 -27480 -2549 -22920
rect 2011 -27480 2035 -22920
rect -2573 -27504 2035 -27480
rect -429 -27936 -109 -27504
rect 2371 -27559 2413 -22841
rect 2649 -27559 2691 -22841
rect 2371 -27881 2691 -27559
rect -2573 -27960 2035 -27936
rect -2573 -32520 -2549 -27960
rect 2011 -32520 2035 -27960
rect -2573 -32544 2035 -32520
rect -429 -32976 -109 -32544
rect 2371 -32599 2413 -27881
rect 2649 -32599 2691 -27881
rect 2371 -32921 2691 -32599
rect -2573 -33000 2035 -32976
rect -2573 -37560 -2549 -33000
rect 2011 -37560 2035 -33000
rect -2573 -37584 2035 -37560
rect -429 -38016 -109 -37584
rect 2371 -37639 2413 -32921
rect 2649 -37639 2691 -32921
rect 2371 -37961 2691 -37639
rect -2573 -38040 2035 -38016
rect -2573 -42600 -2549 -38040
rect 2011 -42600 2035 -38040
rect -2573 -42624 2035 -42600
rect -429 -43056 -109 -42624
rect 2371 -42679 2413 -37961
rect 2649 -42679 2691 -37961
rect 2371 -43001 2691 -42679
rect -2573 -43080 2035 -43056
rect -2573 -47640 -2549 -43080
rect 2011 -47640 2035 -43080
rect -2573 -47664 2035 -47640
rect -429 -48096 -109 -47664
rect 2371 -47719 2413 -43001
rect 2649 -47719 2691 -43001
rect 2371 -48041 2691 -47719
rect -2573 -48120 2035 -48096
rect -2573 -52680 -2549 -48120
rect 2011 -52680 2035 -48120
rect -2573 -52704 2035 -52680
rect -429 -53136 -109 -52704
rect 2371 -52759 2413 -48041
rect 2649 -52759 2691 -48041
rect 2371 -53081 2691 -52759
rect -2573 -53160 2035 -53136
rect -2573 -57720 -2549 -53160
rect 2011 -57720 2035 -53160
rect -2573 -57744 2035 -57720
rect -429 -58176 -109 -57744
rect 2371 -57799 2413 -53081
rect 2649 -57799 2691 -53081
rect 2371 -58121 2691 -57799
rect -2573 -58200 2035 -58176
rect -2573 -62760 -2549 -58200
rect 2011 -62760 2035 -58200
rect -2573 -62784 2035 -62760
rect -429 -63000 -109 -62784
rect 2371 -62839 2413 -58121
rect 2649 -62839 2691 -58121
rect 2371 -63000 2691 -62839
<< properties >>
string FIXED_BBOX -2669 58080 2131 62880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 23.2 l 23.2 val 1.094k carea 2.00 cperi 0.19 nx 1 ny 25 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
