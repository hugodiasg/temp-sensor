** sch_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma_tb-tran.sch
**.subckt sigma_tb-tran
VDD vd GND 1.8
vin in GND 1
V1 clk GND pulse 0 1.8 '0.495/ 10e6 ' '0.01/10e6 ' '0.01/10e6 ' '0.49/10e6 ' '1/10e6 '
x1 gnd_d vpwr clk vd out in vpwr GND sigma-delta
vpwr vpwr GND 1.8
vgndd gnd_d GND 0
C1 out 0 3f m=1
**** begin user architecture code

*cmd step stop
.tran 0.5n 5u
.control
set color0=white
set color1=black
set temp=27
destroy all
run

plot in x1.in_comp x1.out_comp x1.QN
plot clk
plot in
plot out


.endc

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sym # of pins=8
** sym_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/sigma-delta.sch
.subckt sigma-delta  gnd_d vpwr clk vd out in reset_b_dff gnd
*.ipin in
*.iopin gnd
*.iopin clk
*.iopin out
*.iopin reset_b_dff
*.iopin vpwr
*.iopin gnd_d
*.iopin vd
**** begin user architecture code




**** end user architecture code
XC1 in_comp gnd sky130_fd_pr__cap_mim_m3_1 W=27.196 L=27.196 MF=1 m=1
XR2 QN in_comp gnd sky130_fd_pr__res_xhigh_po_0p35 L=37 mult=1 m=1
x2 clk out_comp reset_b_dff gnd_d gnd_d vpwr vpwr out QN sky130_fd_sc_hd__dfrbp_1
XP1 out_comp in_comp vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XN1 out_comp in_comp gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1 in_comp in gnd sky130_fd_pr__res_xhigh_po_0p35 L=37 mult=1 m=1
.ends

.GLOBAL GND
.end
