** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator-pex.sch
**.subckt ask-modulator-pex gnd in out vd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
x1 vd out l0
**** begin user architecture code

* NGSPICE file created from ask-modulator.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN w_n201_n1098# a_n35_500# a_n35_n932#
X0 a_n35_n932# a_n35_500# w_n201_n1098# sky130_fd_pr__res_xhigh_po_0p35 l=5e+06u
C0 a_n35_n932# w_n201_n1098# 1.08fF
C1 a_n35_500# w_n201_n1098# 1.08fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_EZRVX8 m4_n2509_n7390# c2_n2409_n7290# VSUBS
X0 c2_n2409_n7290# m4_n2509_n7390# sky130_fd_pr__cap_mim_m3_2 l=2.33e+07u w=2.33e+07u
X1 c2_n2409_n7290# m4_n2509_n7390# sky130_fd_pr__cap_mim_m3_2 l=2.33e+07u w=2.33e+07u
X2 c2_n2409_n7290# m4_n2509_n7390# sky130_fd_pr__cap_mim_m3_2 l=2.33e+07u w=2.33e+07u
C0 c2_n2409_n7290# m4_n2509_n7390# 108.99fF
C1 c2_n2409_n7290# VSUBS 0.26fF
C2 m4_n2509_n7390# VSUBS 28.74fF
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PWYS4E a_n108_n870# a_n50_n958# w_n278_n1128#  a_50_n870#
X0 a_50_n870# a_n50_n958# a_n108_n870# w_n278_n1128# sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p
+ pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=8.7e+06u l=500000u
C0 a_n108_n870# a_50_n870# 1.03fF
C1 a_50_n870# w_n278_n1128# 0.84fF
C2 a_n108_n870# w_n278_n1128# 0.84fF
C3 a_n50_n958# w_n278_n1128# 0.52fF
.ends

*.subckt ask-modulator in out vd gnd
Xsky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0 gnd vd out sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN
Xsky130_fd_pr__cap_mim_m3_2_EZRVX8_0 out vd gnd sky130_fd_pr__cap_mim_m3_2_EZRVX8
Xsky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5_PWYS4E
*X0 vd.t0 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X1 gnd in.t0 out gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p
*+ ps=1.798e+07u w=0u l=0u
*X2 vd.t2 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X3 vd.t1 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 vd vd.t2 6.883
R1 vd.t1 vd.t0 0.066
R2 vd.t2 vd.t1 0.066
R3 in in.t0 448.598
C0 in out 0.46fF
C1 vd out 7.37fF
C2 in.t0 gnd 0.45fF
C3 vd.t0 gnd 30.94fF
C4 vd.t1 gnd 31.02fF
C5 vd.t2 gnd 173.21fF
C6 out gnd 210.63fF
C7 in gnd 5.53fF
C8 vd gnd 126.57fF
*.ends

**** end user architecture code
**.ends

* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym # of
*+ pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sch
.subckt l0  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.077n m=1
Cs1 p1 net1 10.78f m=1
Cs2 p2 net2 10.54f m=1
Rs1 net1 GND 41.95 m=1
Rs2 net2 GND 5.649 m=1
R1 p2 net3 4.88 m=1
.ends

.GLOBAL GND
.end
