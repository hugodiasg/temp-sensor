magic
tech sky130A
magscale 1 2
timestamp 1668740706
<< nwell >>
rect -683 -969 683 969
<< pmos >>
rect -487 -750 -287 750
rect -229 -750 -29 750
rect 29 -750 229 750
rect 287 -750 487 750
<< pdiff >>
rect -545 738 -487 750
rect -545 -738 -533 738
rect -499 -738 -487 738
rect -545 -750 -487 -738
rect -287 738 -229 750
rect -287 -738 -275 738
rect -241 -738 -229 738
rect -287 -750 -229 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 229 738 287 750
rect 229 -738 241 738
rect 275 -738 287 738
rect 229 -750 287 -738
rect 487 738 545 750
rect 487 -738 499 738
rect 533 -738 545 738
rect 487 -750 545 -738
<< pdiffc >>
rect -533 -738 -499 738
rect -275 -738 -241 738
rect -17 -738 17 738
rect 241 -738 275 738
rect 499 -738 533 738
<< nsubdiff >>
rect -647 899 -551 933
rect 551 899 647 933
rect -647 837 -613 899
rect 613 837 647 899
rect -647 -899 -613 -837
rect 613 -899 647 -837
rect -647 -933 -551 -899
rect 551 -933 647 -899
<< nsubdiffcont >>
rect -551 899 551 933
rect -647 -837 -613 837
rect 613 -837 647 837
rect -551 -933 551 -899
<< poly >>
rect -487 831 -287 847
rect -487 797 -471 831
rect -303 797 -287 831
rect -487 750 -287 797
rect -229 831 -29 847
rect -229 797 -213 831
rect -45 797 -29 831
rect -229 750 -29 797
rect 29 831 229 847
rect 29 797 45 831
rect 213 797 229 831
rect 29 750 229 797
rect 287 831 487 847
rect 287 797 303 831
rect 471 797 487 831
rect 287 750 487 797
rect -487 -797 -287 -750
rect -487 -831 -471 -797
rect -303 -831 -287 -797
rect -487 -847 -287 -831
rect -229 -797 -29 -750
rect -229 -831 -213 -797
rect -45 -831 -29 -797
rect -229 -847 -29 -831
rect 29 -797 229 -750
rect 29 -831 45 -797
rect 213 -831 229 -797
rect 29 -847 229 -831
rect 287 -797 487 -750
rect 287 -831 303 -797
rect 471 -831 487 -797
rect 287 -847 487 -831
<< polycont >>
rect -471 797 -303 831
rect -213 797 -45 831
rect 45 797 213 831
rect 303 797 471 831
rect -471 -831 -303 -797
rect -213 -831 -45 -797
rect 45 -831 213 -797
rect 303 -831 471 -797
<< locali >>
rect -647 899 -551 933
rect 551 899 647 933
rect -647 837 -613 899
rect 613 837 647 899
rect -487 797 -471 831
rect -303 797 -287 831
rect -229 797 -213 831
rect -45 797 -29 831
rect 29 797 45 831
rect 213 797 229 831
rect 287 797 303 831
rect 471 797 487 831
rect -533 738 -499 754
rect -533 -754 -499 -738
rect -275 738 -241 754
rect -275 -754 -241 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 241 738 275 754
rect 241 -754 275 -738
rect 499 738 533 754
rect 499 -754 533 -738
rect -487 -831 -471 -797
rect -303 -831 -287 -797
rect -229 -831 -213 -797
rect -45 -831 -29 -797
rect 29 -831 45 -797
rect 213 -831 229 -797
rect 287 -831 303 -797
rect 471 -831 487 -797
rect -647 -899 -613 -837
rect 613 -899 647 -837
rect -647 -933 -551 -899
rect 551 -933 647 -899
<< viali >>
rect -471 797 -303 831
rect -213 797 -45 831
rect 45 797 213 831
rect 303 797 471 831
rect -533 131 -499 721
rect -275 -295 -241 295
rect -17 131 17 721
rect 241 -295 275 295
rect 499 131 533 721
rect -471 -831 -303 -797
rect -213 -831 -45 -797
rect 45 -831 213 -797
rect 303 -831 471 -797
<< metal1 >>
rect -483 831 -291 837
rect -483 797 -471 831
rect -303 797 -291 831
rect -483 791 -291 797
rect -225 831 -33 837
rect -225 797 -213 831
rect -45 797 -33 831
rect -225 791 -33 797
rect 33 831 225 837
rect 33 797 45 831
rect 213 797 225 831
rect 33 791 225 797
rect 291 831 483 837
rect 291 797 303 831
rect 471 797 483 831
rect 291 791 483 797
rect -539 721 -493 733
rect -539 131 -533 721
rect -499 131 -493 721
rect -23 721 23 733
rect -539 119 -493 131
rect -281 295 -235 307
rect -281 -295 -275 295
rect -241 -295 -235 295
rect -23 131 -17 721
rect 17 131 23 721
rect 493 721 539 733
rect -23 119 23 131
rect 235 295 281 307
rect -281 -307 -235 -295
rect 235 -295 241 295
rect 275 -295 281 295
rect 493 131 499 721
rect 533 131 539 721
rect 493 119 539 131
rect 235 -307 281 -295
rect -483 -797 -291 -791
rect -483 -831 -471 -797
rect -303 -831 -291 -797
rect -483 -837 -291 -831
rect -225 -797 -33 -791
rect -225 -831 -213 -797
rect -45 -831 -33 -797
rect -225 -837 -33 -831
rect 33 -797 225 -791
rect 33 -831 45 -797
rect 213 -831 225 -797
rect 33 -837 225 -831
rect 291 -797 483 -791
rect 291 -831 303 -797
rect 471 -831 483 -797
rect 291 -837 483 -831
<< properties >>
string FIXED_BBOX -630 -916 630 916
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.5 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
