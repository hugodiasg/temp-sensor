magic
tech sky130A
magscale 1 2
timestamp 1645148224
<< error_p >>
rect -2923 -2764 -2863 2764
rect -2843 -2764 -2783 2764
rect 2783 -2764 2843 2764
rect 2863 -2764 2923 2764
<< metal4 >>
rect -8549 2723 -2863 2764
rect -8549 -2723 -3119 2723
rect -2883 -2723 -2863 2723
rect -8549 -2764 -2863 -2723
rect -2843 2723 2843 2764
rect -2843 -2723 2587 2723
rect 2823 -2723 2843 2723
rect -2843 -2764 2843 -2723
rect 2863 2723 8549 2764
rect 2863 -2723 8293 2723
rect 8529 -2723 8549 2723
rect 2863 -2764 8549 -2723
<< via4 >>
rect -3119 -2723 -2883 2723
rect 2587 -2723 2823 2723
rect 8293 -2723 8529 2723
<< mimcap2 >>
rect -8449 2624 -3121 2664
rect -8449 -2624 -7884 2624
rect -3686 -2624 -3121 2624
rect -8449 -2664 -3121 -2624
rect -2743 2624 2585 2664
rect -2743 -2624 -2178 2624
rect 2020 -2624 2585 2624
rect -2743 -2664 2585 -2624
rect 2963 2624 8291 2664
rect 2963 -2624 3528 2624
rect 7726 -2624 8291 2624
rect 2963 -2664 8291 -2624
<< mimcap2contact >>
rect -7884 -2624 -3686 2624
rect -2178 -2624 2020 2624
rect 3528 -2624 7726 2624
<< metal5 >>
rect -3161 2723 -2841 2765
rect -7908 2624 -3662 2648
rect -7908 -2624 -7884 2624
rect -3686 -2624 -3662 2624
rect -7908 -2648 -3662 -2624
rect -3161 -2723 -3119 2723
rect -2883 -2723 -2841 2723
rect 2545 2723 2865 2765
rect -2202 2624 2044 2648
rect -2202 -2624 -2178 2624
rect 2020 -2624 2044 2624
rect -2202 -2648 2044 -2624
rect -3161 -2765 -2841 -2723
rect 2545 -2723 2587 2723
rect 2823 -2723 2865 2723
rect 8251 2723 8571 2765
rect 3504 2624 7750 2648
rect 3504 -2624 3528 2624
rect 7726 -2624 7750 2624
rect 3504 -2648 7750 -2624
rect 2545 -2765 2865 -2723
rect 8251 -2723 8293 2723
rect 8529 -2723 8571 2723
rect 8251 -2765 8571 -2723
<< properties >>
string FIXED_BBOX 2863 -2764 8391 2764
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 26.643 l 26.643 val 1.439k carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
