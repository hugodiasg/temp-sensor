magic
tech sky130A
magscale 1 2
timestamp 1643995581
<< metal1 >>
rect -9000 14200 -3600 14400
rect -9000 13200 -8800 14200
rect -7200 13200 -3600 14200
rect -3000 14200 1800 14400
rect -3000 13200 0 14200
rect 1600 13200 1800 14200
rect -9000 13000 -7000 13200
rect -4800 11520 -4400 13200
rect -3960 12520 -2680 13080
rect -3740 12100 -2680 12520
rect -3180 11920 -2680 12100
rect -3620 11720 -2680 11920
rect -4800 11280 -3420 11520
rect -4800 6900 -4400 11280
rect -3600 6900 -3300 11040
rect -3040 6900 -2680 11720
rect -1720 6900 -1320 13200
rect -200 13000 1800 13200
rect -4700 6700 -4500 6900
rect -3560 6700 -3360 6900
rect -2960 6700 -2760 6900
rect -1660 6700 -1460 6900
<< via1 >>
rect -8800 13200 -7200 14200
rect 0 13200 1600 14200
<< metal2 >>
rect -9000 14200 -7000 14400
rect -9000 13200 -8800 14200
rect -7200 13200 -7000 14200
rect -9000 13000 -7000 13200
rect -200 14200 1800 14400
rect -200 13200 0 14200
rect 1600 13200 1800 14200
rect -200 13000 1800 13200
<< via2 >>
rect -8800 13200 -7200 14200
rect 0 13200 1600 14200
<< metal3 >>
rect -9000 14200 -7000 14400
rect -9000 13200 -8800 14200
rect -7200 13200 -7000 14200
rect -9000 13000 -7000 13200
rect -200 14200 1800 14400
rect -200 13200 0 14200
rect 1600 13200 1800 14200
rect -200 13000 1800 13200
<< via3 >>
rect -8800 13200 -7200 14200
rect 0 13200 1600 14200
<< metal4 >>
rect -9000 29200 -5000 33600
rect -9000 27200 -7000 29200
rect -9000 22800 -4600 27200
rect -9000 20800 -7000 22800
rect -9000 16400 -4400 20800
rect -9000 14200 -7000 16400
rect -9000 13200 -8800 14200
rect -7200 13200 -7000 14200
rect -9000 9600 -7000 13200
rect -200 14200 1800 14400
rect -200 13200 0 14200
rect 1600 13200 1800 14200
rect -200 13000 1800 13200
rect -9000 7600 17000 9600
<< via4 >>
rect 0 13200 1600 14200
<< metal5 >>
rect -1400 31400 2800 33400
rect -1400 29000 1800 31400
rect -200 27400 1800 29000
rect -1200 22600 1800 27400
rect -200 21000 1800 22600
rect -1400 16200 1800 21000
rect -200 14200 1800 16200
rect -200 13200 0 14200
rect 1600 13200 1800 14200
rect -200 13000 1800 13200
use l0  l0_0
timestamp 1643995138
transform 1 0 2300 0 1 10800
box 0 -2000 22600 22600
use sky130_fd_pr__res_high_po_5p73_2BGFUD  XR1
timestamp 1643981260
transform 0 1 -3352 -1 0 13739
box -739 -648 739 648
use sky130_fd_pr__nfet_g5v0d10v5_JF8TZN  XM2
timestamp 1643981260
transform 1 0 -3443 0 1 11493
box -357 -693 357 693
use sky130_fd_pr__cap_mim_m3_2_5KDT2C  XC3
timestamp 1643981260
transform 0 1 -3249 -1 0 18223
box -2801 -2551 2823 2551
use sky130_fd_pr__cap_mim_m3_2_5KDT2C  XC2
timestamp 1643981260
transform 0 1 -3249 -1 0 24623
box -2801 -2551 2823 2551
use sky130_fd_pr__cap_mim_m3_2_5KDT2C  XC1
timestamp 1643981260
transform 0 1 -3249 -1 0 31023
box -2801 -2551 2823 2551
<< labels >>
flabel metal1 -2960 6700 -2760 6900 0 FreeSans 128 0 0 0 gnd
port 0 nsew
flabel metal1 -3560 6700 -3360 6900 0 FreeSans 128 0 0 0 in
port 1 nsew
flabel metal1 -4700 6700 -4500 6900 0 FreeSans 128 0 0 0 out
port 2 nsew
flabel metal1 -1660 6700 -1460 6900 0 FreeSans 128 0 0 0 vd
port 3 nsew
<< properties >>
string l0_0 l0_0
string l0 device
<< end >>
