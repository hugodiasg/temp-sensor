magic
tech sky130A
timestamp 1645758648
<< metal4 >>
rect 209050 265169 265350 265400
rect 209050 264331 257931 265169
rect 258769 264331 259531 265169
rect 260369 264331 261131 265169
rect 261969 264331 262731 265169
rect 263569 264331 264331 265169
rect 265169 264331 265350 265169
rect 209050 263569 265350 264331
rect 209050 262731 257931 263569
rect 258769 262731 259531 263569
rect 260369 262731 261131 263569
rect 261969 262731 262731 263569
rect 263569 262731 264331 263569
rect 265169 262731 265350 263569
rect 209050 261969 265350 262731
rect 209050 261131 257931 261969
rect 258769 261131 259531 261969
rect 260369 261131 261131 261969
rect 261969 261131 262731 261969
rect 263569 261131 264331 261969
rect 265169 261131 265350 261969
rect 209050 260369 265350 261131
rect 209050 259531 257931 260369
rect 258769 259531 259531 260369
rect 260369 259531 261131 260369
rect 261969 259531 262731 260369
rect 263569 259531 264331 260369
rect 265169 259531 265350 260369
rect 209050 258769 265350 259531
rect 209050 257931 257931 258769
rect 258769 257931 259531 258769
rect 260369 257931 261131 258769
rect 261969 257931 262731 258769
rect 263569 257931 264331 258769
rect 265169 257931 265350 258769
rect 209050 257700 265350 257931
<< via4 >>
rect 257931 264331 258769 265169
rect 259531 264331 260369 265169
rect 261131 264331 261969 265169
rect 262731 264331 263569 265169
rect 264331 264331 265169 265169
rect 257931 262731 258769 263569
rect 259531 262731 260369 263569
rect 261131 262731 261969 263569
rect 262731 262731 263569 263569
rect 264331 262731 265169 263569
rect 257931 261131 258769 261969
rect 259531 261131 260369 261969
rect 261131 261131 261969 261969
rect 262731 261131 263569 261969
rect 264331 261131 265169 261969
rect 257931 259531 258769 260369
rect 259531 259531 260369 260369
rect 261131 259531 261969 260369
rect 262731 259531 263569 260369
rect 264331 259531 265169 260369
rect 257931 257931 258769 258769
rect 259531 257931 260369 258769
rect 261131 257931 261969 258769
rect 262731 257931 263569 258769
rect 264331 257931 265169 258769
<< metal5 >>
rect 216000 288300 296000 296000
rect 216000 278100 285800 285800
rect 216000 223699 223699 278100
rect 226199 267900 275600 275600
rect 226199 233899 233899 267900
rect 236399 265169 265400 265400
rect 236399 264331 257931 265169
rect 258769 264331 259531 265169
rect 260369 264331 261131 265169
rect 261969 264331 262731 265169
rect 263569 264331 264331 265169
rect 265169 264331 265400 265169
rect 236399 263569 265400 264331
rect 236399 262731 257931 263569
rect 258769 262731 259531 263569
rect 260369 262731 261131 263569
rect 261969 262731 262731 263569
rect 263569 262731 264331 263569
rect 265169 262731 265400 263569
rect 236399 261969 265400 262731
rect 236399 261131 257931 261969
rect 258769 261131 259531 261969
rect 260369 261131 261131 261969
rect 261969 261131 262731 261969
rect 263569 261131 264331 261969
rect 265169 261131 265400 261969
rect 236399 260369 265400 261131
rect 236399 259531 257931 260369
rect 258769 259531 259531 260369
rect 260369 259531 261131 260369
rect 261969 259531 262731 260369
rect 263569 259531 264331 260369
rect 265169 259531 265400 260369
rect 236399 258769 265400 259531
rect 236399 257931 257931 258769
rect 258769 257931 259531 258769
rect 260369 257931 261131 258769
rect 261969 257931 262731 258769
rect 263569 257931 264331 258769
rect 265169 257931 265400 258769
rect 236399 257700 265400 257931
rect 236399 244099 244099 257700
rect 267900 244099 275600 267900
rect 236399 236399 275600 244099
rect 278100 233899 285800 278100
rect 226199 226199 285800 233899
rect 288300 223699 296000 288300
rect 216000 216000 296000 223699
<< end >>
