** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator-pex_tb-ac.sch
**.subckt ask-modulator-pex_tb-ac
Vdd vd GND DC 3.3 AC 0
Vin net1 GND DC 1.8 AC 1
Vin1 net2 GND DC 1.8 AC 1
R1 ns_in1 net1 50 m=1
R3 ns_out1 GND 50 m=1
R4 ns_out2 net2 50 m=1
R5 ns_in2 GND 50 m=1
x1 vd ns_out1 ns_in1 GND ask-modulator-pex
x2 vd ns_out2 ns_in2 GND ask-modulator-pex
**** begin user architecture code



.ac lin 1MEG 2G 4G
.control
destroy all
set units=degrees
run

set color0=white
set color1=black

let z0=50

* Find two S parameters from test circuit
let s_in1 = v(ns_in1)
let s_out1 = v(ns_out1)
let s_in2 = v(ns_in2)
let s_out2 = v(ns_out2)

* Extract Y parameters
*let StoYDelS = ((1+s_in1)*(1+s_out2)-s_out1*s_in2)*z0
*let y_in1 = ((1+s_out2)*(1-s_in1)+s_out1*s_in2/StoYDelS
*let y_out1=-2*s_out1/StoYDelS
*let y_in2=-2*s_in2/StoYDelS
*let y_out2 = ((1+s_in1)*(1-s_out2)+s_out1+s_in2)/StoYDelS

* Extract Z parameters
let StoZDelS = ((1-s_in1)*(1-s_out2)-s_out1*s_in2)/z0
let z_in1 = ((1+s_in1)*(1-s_out2)+s_out1*s_in2)/StoZDelS
let z_out1 = 2*s_out1/StoZDelS
let z_in2 = 2*s_in2/StoZDelS
let z_out2=((1-s_in1)*(1+s_out2)+s_out1*s_in2)/StoZDelS

*plot z_in1
*plot z_out1
*plot z_in2
plot z_out2 xlimit 2.4G 2.5G
plot ph(z_out2) xlimit 2.4G 2.5G
plot z_out2
plot ph(z_out2)
*plot smith z_out2

.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator-pex.sym # of pins=4
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator-pex.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator-pex.sch
.subckt ask-modulator-pex  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
x1 vd out l0
**** begin user architecture code

* NGSPICE file created from ask-modulator.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN w_n201_n1098# a_n35_500# a_n35_n932#
X0 a_n35_n932# a_n35_500# w_n201_n1098# sky130_fd_pr__res_xhigh_po_0p35 l=5e+06u
C0 a_n35_n932# w_n201_n1098# 1.08fF
C1 a_n35_500# w_n201_n1098# 1.08fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_9XH3MC c2_n2414_n7305# m4_n2514_n7405# VSUBS
X0 c2_n2414_n7305# m4_n2514_n7405# sky130_fd_pr__cap_mim_m3_2 l=2.335e+07u w=2.335e+07u
X1 c2_n2414_n7305# m4_n2514_n7405# sky130_fd_pr__cap_mim_m3_2 l=2.335e+07u w=2.335e+07u
X2 c2_n2414_n7305# m4_n2514_n7405# sky130_fd_pr__cap_mim_m3_2 l=2.335e+07u w=2.335e+07u
C0 m4_n2514_n7405# c2_n2414_n7305# 109.41fF
C1 c2_n2414_n7305# VSUBS 0.26fF
C2 m4_n2514_n7405# VSUBS 28.83fF
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PWYS4E a_n108_n870# a_n50_n958# w_n278_n1128#  a_50_n870#
X0 a_50_n870# a_n50_n958# a_n108_n870# w_n278_n1128# sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p
+ pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=8.7e+06u l=500000u
C0 a_50_n870# a_n108_n870# 1.03fF
C1 a_50_n870# w_n278_n1128# 0.84fF
C2 a_n108_n870# w_n278_n1128# 0.84fF
C3 a_n50_n958# w_n278_n1128# 0.52fF
.ends

*.subckt ask-modulator in out vd gnd
Xsky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0 gnd vd out sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN
Xsky130_fd_pr__cap_mim_m3_2_9XH3MC_0 vd out gnd sky130_fd_pr__cap_mim_m3_2_9XH3MC
Xsky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5_PWYS4E
*X0 vd.t1 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X1 vd.t2 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X2 vd.t0 out sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X3 gnd in.t0 out gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p
*+ ps=1.798e+07u w=0u l=0u
R0 vd vd.t1 6.882
R1 vd.t0 vd.t2 0.066
R2 vd.t1 vd.t0 0.066
R3 in in.t0 448.598
C0 in out 0.46fF
C1 out vd 7.37fF
C2 in.t0 gnd 0.45fF
C3 vd.t2 gnd 31.07fF
C4 vd.t0 gnd 31.16fF
C5 vd.t1 gnd 173.38fF
C6 out gnd 211.18fF
C7 in gnd 5.53fF
C8 vd gnd 126.55fF
*.ends



**** end user architecture code
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym # of
*+ pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sch
.subckt l0  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.077n m=1
Cs1 p1 net1 10.78f m=1
Cs2 p2 net2 10.54f m=1
Rs1 net1 GND 41.95 m=1
Rs2 net2 GND 5.649 m=1
R1 p2 net3 4.88 m=1
.ends

.GLOBAL GND
.end
