* NGSPICE file created from sigma-delta.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VPWR Q Q_N a_543_47# a_1847_47#
+ VNB VPB a_193_47# a_448_47# a_1283_21# a_761_289# a_1108_47# a_27_47#
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=1.5393e+12p ps=1.452e+07u w=1e+06u l=150000u
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X2 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X3 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X5 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X6 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.2225e+12p pd=1.139e+07u as=0p ps=0u w=420000u l=150000u
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_1283_21# a_193_47# 0.04fF
C1 a_761_289# a_1108_47# 0.05fF
C2 VPB a_1847_47# 0.02fF
C3 a_448_47# a_193_47# 0.04fF
C4 VPB RESET_B 0.06fF
C5 Q_N VGND 0.04fF
C6 a_761_289# a_543_47# 0.15fF
C7 a_1283_21# a_1108_47# 0.20fF
C8 a_761_289# VGND 0.06fF
C9 D VGND 0.05fF
C10 a_1283_21# VGND 0.19fF
C11 VPWR Q_N 0.05fF
C12 Q VGND 0.07fF
C13 a_448_47# a_543_47# 0.04fF
C14 a_27_47# RESET_B 0.33fF
C15 a_761_289# VPWR 0.08fF
C16 a_448_47# VGND 0.06fF
C17 VPWR D 0.06fF
C18 VPB a_27_47# 0.09fF
C19 a_1283_21# VPWR 0.12fF
C20 VPWR Q 0.06fF
C21 a_1108_47# a_193_47# 0.10fF
C22 a_543_47# a_193_47# 0.16fF
C23 a_448_47# VPWR 0.05fF
C24 VGND a_193_47# 0.05fF
C25 Q_N a_1847_47# 0.03fF
C26 VPWR a_193_47# 0.40fF
C27 a_1108_47# VGND 0.11fF
C28 a_761_289# RESET_B 0.13fF
C29 a_543_47# VGND 0.10fF
C30 VPB a_761_289# 0.03fF
C31 a_1283_21# a_1847_47# 0.07fF
C32 Q a_1847_47# 0.12fF
C33 a_1283_21# RESET_B 0.23fF
C34 VPB D 0.04fF
C35 VPB a_1283_21# 0.10fF
C36 VPB Q 0.01fF
C37 VPWR a_1108_47# 0.14fF
C38 a_651_413# a_761_289# 0.09fF
C39 VPWR a_543_47# 0.08fF
C40 VPWR VGND 0.12fF
C41 a_761_289# a_27_47# 0.04fF
C42 a_27_47# D 0.09fF
C43 a_1283_21# a_27_47# 0.04fF
C44 RESET_B a_193_47# 0.02fF
C45 VPB CLK 0.02fF
C46 VPB a_193_47# 0.07fF
C47 a_448_47# a_27_47# 0.07fF
C48 a_651_413# a_193_47# 0.01fF
C49 RESET_B a_1108_47# 0.17fF
C50 RESET_B a_543_47# 0.15fF
C51 VPB a_1108_47# 0.04fF
C52 VPB a_543_47# 0.04fF
C53 a_27_47# CLK 0.19fF
C54 a_1847_47# VGND 0.07fF
C55 RESET_B VGND 0.29fF
C56 a_27_47# a_193_47# 0.72fF
C57 VPB VGND 0.07fF
C58 a_651_413# a_543_47# 0.05fF
C59 VPWR a_1847_47# 0.13fF
C60 VPWR RESET_B 0.06fF
C61 a_27_47# a_1108_47# 0.09fF
C62 a_1283_21# Q 0.07fF
C63 a_27_47# a_543_47# 0.05fF
C64 VPB VPWR 0.22fF
C65 a_448_47# D 0.12fF
C66 a_27_47# VGND 0.23fF
C67 a_651_413# VPWR 0.11fF
C68 a_761_289# a_193_47# 0.12fF
C69 D a_193_47# 0.15fF
C70 a_27_47# VPWR 0.12fF
C71 Q_N VNB 0.09fF
C72 VGND VNB 1.18fF
C73 VPWR VNB 1.04fF
C74 RESET_B VNB 0.23fF
C75 D VNB 0.14fF
C76 CLK VNB 0.20fF
C77 VPB VNB 2.11fF
C78 a_448_47# VNB 0.01fF
C79 a_1847_47# VNB 0.14fF
C80 a_1108_47# VNB 0.13fF
C81 a_1283_21# VNB 0.46fF
C82 a_543_47# VNB 0.14fF
C83 a_761_289# VNB 0.11fF
C84 a_193_47# VNB 0.24fF
C85 a_27_47# VNB 0.41fF
.ends

.subckt sky130_fd_pr__pfet_01v8_EFDHR4 a_n33_n397# a_n73_n300# a_15_n300# w_n211_n519#
+ VSUBS
X0 a_15_n300# a_n33_n397# a_n73_n300# w_n211_n519# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
C0 a_15_n300# a_n73_n300# 0.48fF
C1 w_n211_n519# a_n33_n397# 0.18fF
C2 w_n211_n519# a_n73_n300# 0.40fF
C3 w_n211_n519# a_15_n300# 0.13fF
C4 a_n33_n397# a_n73_n300# 0.02fF
C5 a_15_n300# a_n33_n397# 0.02fF
C6 a_15_n300# VSUBS 0.11fF
C7 a_n73_n300# VSUBS 0.02fF
C8 a_n33_n397# VSUBS 0.17fF
C9 w_n211_n519# VSUBS 2.09fF
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_EK42PW a_380_n1032# a_48_600# a_380_600# a_n450_n1032#
+ a_214_n1032# a_214_600# a_48_n1032# a_n284_600# a_n118_600# a_n580_n1162# a_n284_n1032#
+ a_n450_600# a_n118_n1032#
X0 a_380_n1032# a_380_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X1 a_214_n1032# a_214_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X2 a_n284_n1032# a_n284_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X3 a_n450_n1032# a_n450_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X4 a_48_n1032# a_48_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X5 a_n118_n1032# a_n118_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
C0 a_48_600# a_214_600# 0.29fF
C1 a_214_n1032# a_48_n1032# 0.29fF
C2 a_380_600# a_380_n1032# 0.01fF
C3 a_n284_600# a_n284_n1032# 0.01fF
C4 a_n450_600# a_n450_n1032# 0.01fF
C5 a_n118_n1032# a_n284_n1032# 0.29fF
C6 a_n118_600# a_n284_600# 0.29fF
C7 a_48_600# a_48_n1032# 0.01fF
C8 a_n118_600# a_48_600# 0.29fF
C9 a_214_n1032# a_214_600# 0.01fF
C10 a_n118_n1032# a_48_n1032# 0.29fF
C11 a_n450_n1032# a_n284_n1032# 0.29fF
C12 a_n118_600# a_n118_n1032# 0.01fF
C13 a_380_600# a_214_600# 0.29fF
C14 a_n450_600# a_n284_600# 0.29fF
C15 a_214_n1032# a_380_n1032# 0.29fF
C16 a_380_n1032# a_n580_n1162# 0.48fF
C17 a_380_600# a_n580_n1162# 0.46fF
C18 a_214_n1032# a_n580_n1162# 0.31fF
C19 a_214_600# a_n580_n1162# 0.30fF
C20 a_48_n1032# a_n580_n1162# 0.31fF
C21 a_48_600# a_n580_n1162# 0.29fF
C22 a_n118_n1032# a_n580_n1162# 0.31fF
C23 a_n118_600# a_n580_n1162# 0.29fF
C24 a_n284_n1032# a_n580_n1162# 0.31fF
C25 a_n284_600# a_n580_n1162# 0.30fF
C26 a_n450_n1032# a_n580_n1162# 0.52fF
C27 a_n450_600# a_n580_n1162# 0.50fF
.ends

.subckt sky130_fd_pr__nfet_01v8_X78HBF a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
C0 a_15_n100# a_n73_n100# 0.16fF
C1 a_15_n100# a_n33_n188# 0.02fF
C2 a_n33_n188# a_n73_n100# 0.02fF
C3 a_15_n100# a_n175_n274# 0.09fF
C4 a_n73_n100# a_n175_n274# 0.15fF
C5 a_n33_n188# a_n175_n274# 0.36fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_A4KLY5 c1_n2770_n2720# m3_n2870_n2820# VSUBS
X0 c1_n2770_n2720# m3_n2870_n2820# sky130_fd_pr__cap_mim_m3_1 l=2.72e+07u w=2.72e+07u
C0 m3_n2870_n2820# c1_n2770_n2720# 62.23fF
C1 c1_n2770_n2720# VSUBS 2.65fF
C2 m3_n2870_n2820# VSUBS 15.73fF
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_ARMGAU a_380_n1032# a_48_600# a_380_600# a_n450_n1032#
+ a_214_n1032# a_214_600# a_48_n1032# a_n284_600# a_n118_600# a_n580_n1162# a_n284_n1032#
+ a_n450_600# a_n118_n1032#
X0 a_380_n1032# a_380_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X1 a_214_n1032# a_214_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X2 a_n284_n1032# a_n284_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X3 a_n450_n1032# a_n450_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X4 a_48_n1032# a_48_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
X5 a_n118_n1032# a_n118_600# a_n580_n1162# sky130_fd_pr__res_xhigh_po_0p35 l=6e+06u
C0 a_n284_600# a_n284_n1032# 0.01fF
C1 a_n284_600# a_n118_600# 0.29fF
C2 a_n118_n1032# a_n284_n1032# 0.29fF
C3 a_214_n1032# a_380_n1032# 0.29fF
C4 a_n284_600# a_n450_600# 0.29fF
C5 a_214_600# a_380_600# 0.29fF
C6 a_n118_600# a_n118_n1032# 0.01fF
C7 a_n118_n1032# a_48_n1032# 0.29fF
C8 a_214_n1032# a_214_600# 0.01fF
C9 a_n450_n1032# a_n284_n1032# 0.29fF
C10 a_214_n1032# a_48_n1032# 0.29fF
C11 a_48_600# a_n118_600# 0.29fF
C12 a_n450_n1032# a_n450_600# 0.01fF
C13 a_48_600# a_214_600# 0.29fF
C14 a_380_600# a_380_n1032# 0.01fF
C15 a_48_600# a_48_n1032# 0.01fF
C16 a_380_n1032# a_n580_n1162# 0.48fF
C17 a_380_600# a_n580_n1162# 0.46fF
C18 a_214_n1032# a_n580_n1162# 0.31fF
C19 a_214_600# a_n580_n1162# 0.30fF
C20 a_48_n1032# a_n580_n1162# 0.31fF
C21 a_48_600# a_n580_n1162# 0.29fF
C22 a_n118_n1032# a_n580_n1162# 0.31fF
C23 a_n118_600# a_n580_n1162# 0.29fF
C24 a_n284_n1032# a_n580_n1162# 0.31fF
C25 a_n284_600# a_n580_n1162# 0.30fF
C26 a_n450_n1032# a_n580_n1162# 0.52fF
C27 a_n450_600# a_n580_n1162# 0.50fF
.ends

.subckt sigma-delta in out clk reset_b_dff vd vpwr gnd
Xx1 clk out_comp reset_b_dff gnd vpwr Q out x1/a_543_47# x1/a_1847_47# gnd vpwr x1/a_193_47#
+ x1/a_448_47# x1/a_1283_21# x1/a_761_289# x1/a_1108_47# x1/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_pr__pfet_01v8_EFDHR4_0 in_comp vd out_comp vd gnd sky130_fd_pr__pfet_01v8_EFDHR4
XXR2 Q m1_n1710_5800# m1_n1400_5790# in_comp m1_n1550_4170# m1_n1400_5790# m1_n1550_4170#
+ m1_n2050_5780# m1_n1710_5800# gnd m1_n1890_4160# m1_n2050_5780# m1_n1890_4160# sky130_fd_pr__res_xhigh_po_0p35_EK42PW
XXN1 gnd in_comp out_comp gnd sky130_fd_pr__nfet_01v8_X78HBF
XXC1 in_comp gnd gnd sky130_fd_pr__cap_mim_m3_1_A4KLY5
Xsky130_fd_pr__res_xhigh_po_0p35_ARMGAU_0 in_comp m1_n3250_5800# m1_n2930_5790# in
+ m1_n3070_4170# m1_n2930_5790# m1_n3070_4170# m1_n3590_5800# m1_n3250_5800# gnd m1_n3420_4160#
+ m1_n3590_5800# m1_n3420_4160# sky130_fd_pr__res_xhigh_po_0p35_ARMGAU
X0 in_comp gnd.t0 sky130_fd_pr__cap_mim_m3_1 l=0u w=0u
X1 vpwr clk.t0 x1/a_27_47# vpwr sky130_fd_pr__pfet_01v8_hvt ad=1.5393e+12p pd=1.452e+07u as=1.664e+11p ps=1.8e+06u w=0u l=0u
X2 x1/a_1462_47# reset_b_dff.t1 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=1.5125e+12p ps=1.397e+07u w=0u l=0u
X3 gnd clk.t1 x1/a_27_47# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=0u l=0u
X4 x1/a_1283_21# reset_b_dff.t2 vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=0u l=0u
X5 x1/a_651_413# reset_b_dff.t3 vpwr vpwr sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=0u l=0u
X6 gnd reset_b_dff.t0 x1/a_805_47# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=0u l=0u
R0 vpwr.n4 vpwr 6628.29
R1 vpwr.n3 vpwr.n0 583.1
R2 vpwr.n4 vpwr.n2 375
R3 vpwr.n5 vpwr.n1 264.705
R4 vpwr vpwr.n3 230.841
R5 vpwr.n6 vpwr.n5 213.235
R6 vpwr.n5 vpwr.n4 185
R7 vpwr.n3 vpwr.n2 95
R8 vpwr vpwr 1.66
R9 vpwr.n7 vpwr 0.366
R10 vpwr vpwr.n7 0.033
R11 vpwr.n2 vpwr.n1 0.003
R12 vpwr.n7 vpwr.n6 0.002
R13 vpwr.n1 vpwr.n0 0.002
R14 vpwr.n6 vpwr.n0 0.002
R15 gnd.n6 gnd.n3 568.151
R16 gnd.n17 gnd.n13 568.151
R17 gnd.n20 gnd.n19 442.745
R18 gnd.n10 gnd.n9 442.728
R19 gnd.n35 gnd.n34 71.545
R20 gnd.n32 gnd.n31 71.491
R21 gnd.n40 gnd 5.358
R22 gnd gnd.n40 3.286
R23 gnd.n39 gnd 2.523
R24 gnd.n38 gnd.n37 1.736
R25 gnd.n23 gnd.n22 1.17
R26 gnd.n38 gnd.n23 0.853
R27 gnd.n23 gnd.t0 0.786
R28 gnd.n11 gnd.n1 0.65
R29 gnd.n37 gnd 0.427
R30 gnd.n20 gnd.n11 0.412
R31 gnd.n21 gnd.n20 0.399
R32 gnd.n37 gnd.n36 0.166
R33 gnd.n22 gnd.n21 0.111
R34 gnd.n34 gnd.n33 0.109
R35 gnd.n31 gnd.n30 0.109
R36 gnd.n39 gnd.n38 0.082
R37 gnd.n25 gnd.n24 0.042
R38 gnd.n27 gnd.n26 0.024
R39 gnd.n26 gnd.n25 0.02
R40 gnd.n11 gnd.n10 0.017
R41 gnd.n3 gnd.n2 0.014
R42 gnd.n13 gnd.n12 0.014
R43 gnd.n8 gnd.n7 0.006
R44 gnd.n16 gnd.n15 0.006
R45 gnd.n6 gnd.n5 0.006
R46 gnd.n18 gnd.n17 0.006
R47 gnd.n9 gnd.n8 0.006
R48 gnd.n5 gnd.n4 0.006
R49 gnd.n15 gnd.n14 0.006
R50 gnd.n19 gnd.n18 0.006
R51 gnd.n7 gnd.n6 0.002
R52 gnd.n17 gnd.n16 0.002
R53 gnd.n32 gnd.n29 0.001
R54 gnd.n29 gnd.n28 0.001
R55 gnd.n28 gnd.n27 0.001
R56 gnd.n40 gnd.n39 0.001
R57 gnd.n36 gnd.n35 0.001
R58 gnd.n36 gnd.n32 0.001
R59 gnd.n1 gnd.n0 0.001
R60 reset_b_dff.n4 reset_b_dff.t3 413.312
R61 reset_b_dff.n12 reset_b_dff.t2 344.005
R62 reset_b_dff.n1 reset_b_dff.t1 187.32
R63 reset_b_dff.n13 reset_b_dff.n12 152
R64 reset_b_dff.n4 reset_b_dff.t0 126.126
R65 reset_b_dff.n1 reset_b_dff.n0 73.206
R66 reset_b_dff.n14 reset_b_dff 14.017
R67 reset_b_dff.n5 reset_b_dff.n4 10.648
R68 reset_b_dff.n8 reset_b_dff.n7 9.3
R69 reset_b_dff.n11 reset_b_dff.n10 9.3
R70 reset_b_dff.n12 reset_b_dff.n11 9.3
R71 reset_b_dff.n12 reset_b_dff.n1 9.159
R72 reset_b_dff.n15 reset_b_dff 7.772
R73 reset_b_dff.n9 reset_b_dff.n2 4.65
R74 reset_b_dff.n14 reset_b_dff 4.533
R75 reset_b_dff reset_b_dff.n13 3.113
R76 reset_b_dff.n15 reset_b_dff.n14 3.033
R77 reset_b_dff reset_b_dff.n6 2.366
R78 reset_b_dff.n13 reset_b_dff.n0 1.556
R79 reset_b_dff.n7 reset_b_dff.n2 1.556
R80 reset_b_dff.n11 reset_b_dff.n0 1.383
R81 reset_b_dff.n11 reset_b_dff.n2 1.383
R82 reset_b_dff.n7 reset_b_dff 1.383
R83 reset_b_dff.n6 reset_b_dff 0.58
R84 reset_b_dff.n5 reset_b_dff 0.271
R85 reset_b_dff.n3 reset_b_dff 0.195
R86 reset_b_dff.n6 reset_b_dff.n5 0.082
R87 reset_b_dff.n16 reset_b_dff.n15 0.045
R88 reset_b_dff.n10 reset_b_dff.n3 0.026
R89 reset_b_dff.n8 reset_b_dff 0.025
R90 reset_b_dff.n9 reset_b_dff.n8 0.011
R91 reset_b_dff.n10 reset_b_dff.n9 0.01
R92 reset_b_dff.n16 reset_b_dff 0.008
R93 reset_b_dff.n3 reset_b_dff 0.006
R94 reset_b_dff reset_b_dff.n16 0.005
R95 clk.n0 clk.t0 294.554
R96 clk.n0 clk.t1 211.008
R97 clk.n1 clk.n0 76
R98 clk.n1 clk 10.422
R99 clk.n1 clk 8.987
R100 clk clk.n1 2.011
R101 out out 4.827
C0 x1/a_1283_21# Q 0.02fF
C1 m1_n2930_5790# m1_n1710_5800# 0.02fF
C2 out_comp clk 0.07fF
C3 reset_b_dff out 0.04fF
C4 gnd x1/a_1847_47# 0.02fF
C5 in_comp reset_b_dff 0.02fF
C6 gnd in 0.15fF
C7 gnd m1_n1550_4170# 0.01fF
C8 gnd clk 0.06fF
C9 vd x1/a_1847_47# 0.01fF
C10 out x1/a_761_289# 0.02fF
C11 out Q 0.12fF
C12 out_comp x1/a_543_47# 0.01fF
C13 vd clk 0.03fF
C14 in_comp Q 0.27fF
C15 x1/a_27_47# vpwr 0.03fF
C16 gnd out_comp 0.34fF
C17 x1/a_1108_47# out_comp 0.01fF
C18 gnd m1_n1890_4160# -0.03fF
C19 x1/a_193_47# out 0.04fF
C20 in vpwr 0.02fF
C21 gnd m1_n2050_5780# 0.01fF
C22 vd out_comp 0.70fF
C23 gnd x1/a_1108_47# 0.01fF
C24 clk vpwr 0.07fF
C25 m1_n2050_5780# m1_n3250_5800# 0.02fF
C26 x1/a_27_47# Q 0.01fF
C27 m1_n3420_4160# gnd 0.04fF
C28 vd gnd 0.66fF
C29 gnd m1_n3250_5800# 0.01fF
C30 gnd m1_n1400_5790# 0.03fF
C31 x1/a_1283_21# out 0.03fF
C32 out_comp vpwr 0.10fF
C33 m1_n1550_4170# Q 0.04fF
C34 reset_b_dff out_comp 0.22fF
C35 gnd vpwr 0.16fF
C36 m1_n2930_5790# in_comp 0.01fF
C37 gnd reset_b_dff 0.13fF
C38 reset_b_dff x1/a_1108_47# 0.01fF
C39 gnd m1_n1710_5800# 0.01fF
C40 vd vpwr 0.05fF
C41 x1/a_761_289# out_comp 0.01fF
C42 Q out_comp 0.02fF
C43 m1_n1890_4160# Q 0.03fF
C44 vd reset_b_dff 0.24fF
C45 m1_n1400_5790# m1_n1710_5800# 0.02fF
C46 gnd Q 0.27fF
C47 x1/a_1108_47# Q 0.01fF
C48 x1/a_193_47# out_comp 0.03fF
C49 x1/a_27_47# out 0.08fF
C50 vd Q 0.01fF
C51 reset_b_dff vpwr 0.01fF
C52 x1/a_1847_47# out 0.02fF
C53 in in_comp 0.14fF
C54 x1/a_1283_21# out_comp 0.02fF
C55 out clk 0.14fF
C56 in_comp m1_n1550_4170# 0.12fF
C57 x1/a_448_47# out_comp -0.02fF
C58 Q vpwr 0.18fF
C59 gnd x1/a_1283_21# 0.02fF
C60 reset_b_dff Q 0.02fF
C61 vd x1/a_1283_21# 0.02fF
C62 out out_comp 0.31fF
C63 out x1/a_543_47# 0.02fF
C64 in_comp out_comp 0.43fF
C65 m1_n2930_5790# m1_n2050_5780# 0.06fF
C66 m1_n1890_4160# in_comp 0.18fF
C67 gnd m1_n2930_5790# 0.01fF
C68 in_comp m1_n3070_4170# 0.19fF
C69 x1/a_27_47# clk 0.03fF
C70 in_comp m1_n2050_5780# 0.01fF
C71 gnd out 0.07fF
C72 out x1/a_1108_47# 0.02fF
C73 gnd in_comp 0.78fF
C74 vd out 0.07fF
C75 m1_n3420_4160# in_comp 0.14fF
C76 vd in_comp 0.22fF
C77 x1/a_193_47# Q 0.01fF
C78 x1/a_27_47# out_comp 0.09fF
C79 gnd x1/a_27_47# -0.02fF
C80 out vpwr 0.38fF
C81 in_comp 0 7.34fF
C82 gnd.t0 0 59.96fF
C83 gnd.n0 0 1.56fF $ **FLOATING
C84 gnd.n1 0 0.14fF $ **FLOATING
C85 gnd.n2 0 0.11fF $ **FLOATING
C86 gnd.n3 0 1.53fF $ **FLOATING
C87 gnd.n4 0 0.09fF $ **FLOATING
C88 gnd.n5 0 0.11fF $ **FLOATING
C89 gnd.n6 0 1.30fF $ **FLOATING
C90 gnd.n7 0 1.30fF $ **FLOATING
C91 gnd.n8 0 0.11fF $ **FLOATING
C92 gnd.n9 0 0.09fF $ **FLOATING
C93 gnd.n10 0 0.05fF $ **FLOATING
C94 gnd.n11 0 0.16fF $ **FLOATING
C95 gnd.n12 0 0.11fF $ **FLOATING
C96 gnd.n13 0 1.53fF $ **FLOATING
C97 gnd.n14 0 0.09fF $ **FLOATING
C98 gnd.n15 0 0.11fF $ **FLOATING
C99 gnd.n16 0 1.30fF $ **FLOATING
C100 gnd.n17 0 1.30fF $ **FLOATING
C101 gnd.n18 0 0.11fF $ **FLOATING
C102 gnd.n19 0 0.09fF $ **FLOATING
C103 gnd.n20 0 0.20fF $ **FLOATING
C104 gnd.n21 0 1.66fF $ **FLOATING
C105 gnd.n22 0 0.32fF $ **FLOATING
C106 gnd.n23 0 1.73fF $ **FLOATING
C107 gnd.n24 0 0.03fF $ **FLOATING
C108 gnd.n25 0 0.03fF $ **FLOATING
C109 gnd.n27 0 0.19fF $ **FLOATING
C110 gnd.n28 0 0.03fF $ **FLOATING
C111 gnd.n29 0 0.01fF $ **FLOATING
C112 gnd.n30 0 0.17fF $ **FLOATING
C113 gnd.n31 0 0.02fF $ **FLOATING
C114 gnd.n32 0 0.02fF $ **FLOATING
C115 gnd.n33 0 0.17fF $ **FLOATING
C116 gnd.n34 0 0.02fF $ **FLOATING
C117 gnd.n35 0 0.02fF $ **FLOATING
C118 gnd.n36 0 0.11fF $ **FLOATING
C119 gnd.n37 0 0.56fF $ **FLOATING
C120 gnd.n38 0 0.49fF $ **FLOATING
C121 gnd.n39 0 0.29fF $ **FLOATING
C122 gnd.n40 0 0.24fF $ **FLOATING
C123 vpwr.n0 0 0.04fF $ **FLOATING
C124 vpwr.n2 0 0.03fF $ **FLOATING
C125 vpwr.n3 0 2.03fF $ **FLOATING
C126 vpwr.n4 0 0.06fF $ **FLOATING
C127 vpwr.n6 0 0.03fF $ **FLOATING
C128 vpwr.n7 0 0.93fF $ **FLOATING
C129 m1_n2930_5790# 0 0.75fF
C130 m1_n3070_4170# 0 0.70fF
C131 m1_n3250_5800# 0 0.64fF
C132 m1_n3420_4160# 0 0.65fF
C133 in 0 1.30fF
C134 m1_n3590_5800# 0 0.86fF
C135 m1_n1400_5790# 0 0.81fF
C136 m1_n1550_4170# 0 0.70fF
C137 m1_n1710_5800# 0 0.65fF
C138 m1_n1890_4160# 0 0.74fF
C139 m1_n2050_5780# 0 0.80fF
C140 out_comp 0 2.24fF
C141 vd 0 7.26fF
C142 out 0 0.41fF
C143 Q 0 1.90fF
C144 gnd 0 15.27fF
C145 reset_b_dff 0 1.53fF
C146 clk 0 0.75fF
C147 vpwr 0 4.81fF
C148 x1/a_448_47# 0 0.01fF
C149 x1/a_1847_47# 0 0.14fF
C150 x1/a_1108_47# 0 0.13fF
C151 x1/a_1283_21# 0 0.46fF
C152 x1/a_543_47# 0 0.14fF
C153 x1/a_761_289# 0 0.11fF
C154 x1/a_193_47# 0 0.24fF
C155 x1/a_27_47# 0 0.41fF
.ends

