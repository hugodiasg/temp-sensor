magic
tech sky130A
magscale 1 2
timestamp 1644767790
<< metal4 >>
rect -2589 7589 2589 7630
rect -2589 2651 2333 7589
rect 2569 2651 2589 7589
rect -2589 2610 2589 2651
rect -2589 2469 2589 2510
rect -2589 -2469 2333 2469
rect 2569 -2469 2589 2469
rect -2589 -2510 2589 -2469
rect -2589 -2651 2589 -2610
rect -2589 -7589 2333 -2651
rect 2569 -7589 2589 -2651
rect -2589 -7630 2589 -7589
<< via4 >>
rect 2333 2651 2569 7589
rect 2333 -2469 2569 2469
rect 2333 -7589 2569 -2651
<< mimcap2 >>
rect -2489 7490 2331 7530
rect -2489 2750 -1975 7490
rect 1817 2750 2331 7490
rect -2489 2710 2331 2750
rect -2489 2370 2331 2410
rect -2489 -2370 -1975 2370
rect 1817 -2370 2331 2370
rect -2489 -2410 2331 -2370
rect -2489 -2750 2331 -2710
rect -2489 -7490 -1975 -2750
rect 1817 -7490 2331 -2750
rect -2489 -7530 2331 -7490
<< mimcap2contact >>
rect -1975 2750 1817 7490
rect -1975 -2370 1817 2370
rect -1975 -7490 1817 -2750
<< metal5 >>
rect -239 7514 81 7680
rect 2291 7589 2611 7680
rect -1999 7490 1841 7514
rect -1999 2750 -1975 7490
rect 1817 2750 1841 7490
rect -1999 2726 1841 2750
rect -239 2394 81 2726
rect 2291 2651 2333 7589
rect 2569 2651 2611 7589
rect 2291 2469 2611 2651
rect -1999 2370 1841 2394
rect -1999 -2370 -1975 2370
rect 1817 -2370 1841 2370
rect -1999 -2394 1841 -2370
rect -239 -2726 81 -2394
rect 2291 -2469 2333 2469
rect 2569 -2469 2611 2469
rect 2291 -2651 2611 -2469
rect -1999 -2750 1841 -2726
rect -1999 -7490 -1975 -2750
rect 1817 -7490 1841 -2750
rect -1999 -7514 1841 -7490
rect -239 -7680 81 -7514
rect 2291 -7589 2333 -2651
rect 2569 -7589 2611 -2651
rect 2291 -7680 2611 -7589
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2589 2610 2431 7630
string parameters w 24.1 l 24.1 val 1.179k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
string library sky130
<< end >>
