magic
tech sky130A
magscale 1 2
timestamp 1646425465
<< metal4 >>
rect -2599 7619 2599 7660
rect -2599 2661 2343 7619
rect 2579 2661 2599 7619
rect -2599 2620 2599 2661
rect -2599 2479 2599 2520
rect -2599 -2479 2343 2479
rect 2579 -2479 2599 2479
rect -2599 -2520 2599 -2479
rect -2599 -2661 2599 -2620
rect -2599 -7619 2343 -2661
rect 2579 -7619 2599 -2661
rect -2599 -7660 2599 -7619
<< via4 >>
rect 2343 2661 2579 7619
rect 2343 -2479 2579 2479
rect 2343 -7619 2579 -2661
<< mimcap2 >>
rect -2499 7520 2341 7560
rect -2499 2760 -1983 7520
rect 1825 2760 2341 7520
rect -2499 2720 2341 2760
rect -2499 2380 2341 2420
rect -2499 -2380 -1983 2380
rect 1825 -2380 2341 2380
rect -2499 -2420 2341 -2380
rect -2499 -2760 2341 -2720
rect -2499 -7520 -1983 -2760
rect 1825 -7520 2341 -2760
rect -2499 -7560 2341 -7520
<< mimcap2contact >>
rect -1983 2760 1825 7520
rect -1983 -2380 1825 2380
rect -1983 -7520 1825 -2760
<< metal5 >>
rect -239 7544 81 7710
rect 2301 7619 2621 7710
rect -2007 7520 1849 7544
rect -2007 2760 -1983 7520
rect 1825 2760 1849 7520
rect -2007 2736 1849 2760
rect -239 2404 81 2736
rect 2301 2661 2343 7619
rect 2579 2661 2621 7619
rect 2301 2479 2621 2661
rect -2007 2380 1849 2404
rect -2007 -2380 -1983 2380
rect 1825 -2380 1849 2380
rect -2007 -2404 1849 -2380
rect -239 -2736 81 -2404
rect 2301 -2479 2343 2479
rect 2579 -2479 2621 2479
rect 2301 -2661 2621 -2479
rect -2007 -2760 1849 -2736
rect -2007 -7520 -1983 -2760
rect 1825 -7520 1849 -2760
rect -2007 -7544 1849 -7520
rect -239 -7710 81 -7544
rect 2301 -7619 2343 -2661
rect 2579 -7619 2621 -2661
rect 2301 -7710 2621 -7619
<< properties >>
string FIXED_BBOX -2599 2620 2441 7660
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.2 l 24.2 val 1.189k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
