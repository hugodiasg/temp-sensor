magic
tech sky130A
magscale 1 2
timestamp 1661128600
<< pwell >>
rect -1457 -310 1457 310
<< nmos >>
rect -1261 -100 -1061 100
rect -1003 -100 -803 100
rect -745 -100 -545 100
rect -487 -100 -287 100
rect -229 -100 -29 100
rect 29 -100 229 100
rect 287 -100 487 100
rect 545 -100 745 100
rect 803 -100 1003 100
rect 1061 -100 1261 100
<< ndiff >>
rect -1319 88 -1261 100
rect -1319 -88 -1307 88
rect -1273 -88 -1261 88
rect -1319 -100 -1261 -88
rect -1061 88 -1003 100
rect -1061 -88 -1049 88
rect -1015 -88 -1003 88
rect -1061 -100 -1003 -88
rect -803 88 -745 100
rect -803 -88 -791 88
rect -757 -88 -745 88
rect -803 -100 -745 -88
rect -545 88 -487 100
rect -545 -88 -533 88
rect -499 -88 -487 88
rect -545 -100 -487 -88
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
rect 487 88 545 100
rect 487 -88 499 88
rect 533 -88 545 88
rect 487 -100 545 -88
rect 745 88 803 100
rect 745 -88 757 88
rect 791 -88 803 88
rect 745 -100 803 -88
rect 1003 88 1061 100
rect 1003 -88 1015 88
rect 1049 -88 1061 88
rect 1003 -100 1061 -88
rect 1261 88 1319 100
rect 1261 -88 1273 88
rect 1307 -88 1319 88
rect 1261 -100 1319 -88
<< ndiffc >>
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
<< psubdiff >>
rect -1421 240 -1325 274
rect 1325 240 1421 274
rect -1421 178 -1387 240
rect 1387 178 1421 240
rect -1421 -240 -1387 -178
rect 1387 -240 1421 -178
rect -1421 -274 -1325 -240
rect 1325 -274 1421 -240
<< psubdiffcont >>
rect -1325 240 1325 274
rect -1421 -178 -1387 178
rect 1387 -178 1421 178
rect -1325 -274 1325 -240
<< poly >>
rect -1261 172 -1061 188
rect -1261 138 -1245 172
rect -1077 138 -1061 172
rect -1261 100 -1061 138
rect -1003 172 -803 188
rect -1003 138 -987 172
rect -819 138 -803 172
rect -1003 100 -803 138
rect -745 172 -545 188
rect -745 138 -729 172
rect -561 138 -545 172
rect -745 100 -545 138
rect -487 172 -287 188
rect -487 138 -471 172
rect -303 138 -287 172
rect -487 100 -287 138
rect -229 172 -29 188
rect -229 138 -213 172
rect -45 138 -29 172
rect -229 100 -29 138
rect 29 172 229 188
rect 29 138 45 172
rect 213 138 229 172
rect 29 100 229 138
rect 287 172 487 188
rect 287 138 303 172
rect 471 138 487 172
rect 287 100 487 138
rect 545 172 745 188
rect 545 138 561 172
rect 729 138 745 172
rect 545 100 745 138
rect 803 172 1003 188
rect 803 138 819 172
rect 987 138 1003 172
rect 803 100 1003 138
rect 1061 172 1261 188
rect 1061 138 1077 172
rect 1245 138 1261 172
rect 1061 100 1261 138
rect -1261 -138 -1061 -100
rect -1261 -172 -1245 -138
rect -1077 -172 -1061 -138
rect -1261 -188 -1061 -172
rect -1003 -138 -803 -100
rect -1003 -172 -987 -138
rect -819 -172 -803 -138
rect -1003 -188 -803 -172
rect -745 -138 -545 -100
rect -745 -172 -729 -138
rect -561 -172 -545 -138
rect -745 -188 -545 -172
rect -487 -138 -287 -100
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -487 -188 -287 -172
rect -229 -138 -29 -100
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect -229 -188 -29 -172
rect 29 -138 229 -100
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 29 -188 229 -172
rect 287 -138 487 -100
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 287 -188 487 -172
rect 545 -138 745 -100
rect 545 -172 561 -138
rect 729 -172 745 -138
rect 545 -188 745 -172
rect 803 -138 1003 -100
rect 803 -172 819 -138
rect 987 -172 1003 -138
rect 803 -188 1003 -172
rect 1061 -138 1261 -100
rect 1061 -172 1077 -138
rect 1245 -172 1261 -138
rect 1061 -188 1261 -172
<< polycont >>
rect -1245 138 -1077 172
rect -987 138 -819 172
rect -729 138 -561 172
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect 561 138 729 172
rect 819 138 987 172
rect 1077 138 1245 172
rect -1245 -172 -1077 -138
rect -987 -172 -819 -138
rect -729 -172 -561 -138
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
rect 561 -172 729 -138
rect 819 -172 987 -138
rect 1077 -172 1245 -138
<< locali >>
rect -1421 240 -1325 274
rect 1325 240 1421 274
rect -1421 178 -1387 240
rect 1387 178 1421 240
rect -1261 138 -1245 172
rect -1077 138 -1061 172
rect -1003 138 -987 172
rect -819 138 -803 172
rect -745 138 -729 172
rect -561 138 -545 172
rect -487 138 -471 172
rect -303 138 -287 172
rect -229 138 -213 172
rect -45 138 -29 172
rect 29 138 45 172
rect 213 138 229 172
rect 287 138 303 172
rect 471 138 487 172
rect 545 138 561 172
rect 729 138 745 172
rect 803 138 819 172
rect 987 138 1003 172
rect 1061 138 1077 172
rect 1245 138 1261 172
rect -1307 88 -1273 104
rect -1307 -104 -1273 -88
rect -1049 88 -1015 104
rect -1049 -104 -1015 -88
rect -791 88 -757 104
rect -791 -104 -757 -88
rect -533 88 -499 104
rect -533 -104 -499 -88
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect 499 88 533 104
rect 499 -104 533 -88
rect 757 88 791 104
rect 757 -104 791 -88
rect 1015 88 1049 104
rect 1015 -104 1049 -88
rect 1273 88 1307 104
rect 1273 -104 1307 -88
rect -1261 -172 -1245 -138
rect -1077 -172 -1061 -138
rect -1003 -172 -987 -138
rect -819 -172 -803 -138
rect -745 -172 -729 -138
rect -561 -172 -545 -138
rect -487 -172 -471 -138
rect -303 -172 -287 -138
rect -229 -172 -213 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 213 -172 229 -138
rect 287 -172 303 -138
rect 471 -172 487 -138
rect 545 -172 561 -138
rect 729 -172 745 -138
rect 803 -172 819 -138
rect 987 -172 1003 -138
rect 1061 -172 1077 -138
rect 1245 -172 1261 -138
rect -1421 -240 -1387 -178
rect 1387 -240 1421 -178
rect -1421 -274 -1325 -240
rect 1325 -274 1421 -240
<< viali >>
rect -1245 138 -1077 172
rect -987 138 -819 172
rect -729 138 -561 172
rect -471 138 -303 172
rect -213 138 -45 172
rect 45 138 213 172
rect 303 138 471 172
rect 561 138 729 172
rect 819 138 987 172
rect 1077 138 1245 172
rect -1307 -88 -1273 88
rect -1049 -88 -1015 88
rect -791 -88 -757 88
rect -533 -88 -499 88
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect 499 -88 533 88
rect 757 -88 791 88
rect 1015 -88 1049 88
rect 1273 -88 1307 88
rect -1245 -172 -1077 -138
rect -987 -172 -819 -138
rect -729 -172 -561 -138
rect -471 -172 -303 -138
rect -213 -172 -45 -138
rect 45 -172 213 -138
rect 303 -172 471 -138
rect 561 -172 729 -138
rect 819 -172 987 -138
rect 1077 -172 1245 -138
<< metal1 >>
rect -1257 172 -1065 178
rect -1257 138 -1245 172
rect -1077 138 -1065 172
rect -1257 132 -1065 138
rect -999 172 -807 178
rect -999 138 -987 172
rect -819 138 -807 172
rect -999 132 -807 138
rect -741 172 -549 178
rect -741 138 -729 172
rect -561 138 -549 172
rect -741 132 -549 138
rect -483 172 -291 178
rect -483 138 -471 172
rect -303 138 -291 172
rect -483 132 -291 138
rect -225 172 -33 178
rect -225 138 -213 172
rect -45 138 -33 172
rect -225 132 -33 138
rect 33 172 225 178
rect 33 138 45 172
rect 213 138 225 172
rect 33 132 225 138
rect 291 172 483 178
rect 291 138 303 172
rect 471 138 483 172
rect 291 132 483 138
rect 549 172 741 178
rect 549 138 561 172
rect 729 138 741 172
rect 549 132 741 138
rect 807 172 999 178
rect 807 138 819 172
rect 987 138 999 172
rect 807 132 999 138
rect 1065 172 1257 178
rect 1065 138 1077 172
rect 1245 138 1257 172
rect 1065 132 1257 138
rect -1313 88 -1267 100
rect -1313 -88 -1307 88
rect -1273 -88 -1267 88
rect -1313 -100 -1267 -88
rect -1055 88 -1009 100
rect -1055 -88 -1049 88
rect -1015 -88 -1009 88
rect -1055 -100 -1009 -88
rect -797 88 -751 100
rect -797 -88 -791 88
rect -757 -88 -751 88
rect -797 -100 -751 -88
rect -539 88 -493 100
rect -539 -88 -533 88
rect -499 -88 -493 88
rect -539 -100 -493 -88
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect 493 88 539 100
rect 493 -88 499 88
rect 533 -88 539 88
rect 493 -100 539 -88
rect 751 88 797 100
rect 751 -88 757 88
rect 791 -88 797 88
rect 751 -100 797 -88
rect 1009 88 1055 100
rect 1009 -88 1015 88
rect 1049 -88 1055 88
rect 1009 -100 1055 -88
rect 1267 88 1313 100
rect 1267 -88 1273 88
rect 1307 -88 1313 88
rect 1267 -100 1313 -88
rect -1257 -138 -1065 -132
rect -1257 -172 -1245 -138
rect -1077 -172 -1065 -138
rect -1257 -178 -1065 -172
rect -999 -138 -807 -132
rect -999 -172 -987 -138
rect -819 -172 -807 -138
rect -999 -178 -807 -172
rect -741 -138 -549 -132
rect -741 -172 -729 -138
rect -561 -172 -549 -138
rect -741 -178 -549 -172
rect -483 -138 -291 -132
rect -483 -172 -471 -138
rect -303 -172 -291 -138
rect -483 -178 -291 -172
rect -225 -138 -33 -132
rect -225 -172 -213 -138
rect -45 -172 -33 -138
rect -225 -178 -33 -172
rect 33 -138 225 -132
rect 33 -172 45 -138
rect 213 -172 225 -138
rect 33 -178 225 -172
rect 291 -138 483 -132
rect 291 -172 303 -138
rect 471 -172 483 -138
rect 291 -178 483 -172
rect 549 -138 741 -132
rect 549 -172 561 -138
rect 729 -172 741 -138
rect 549 -178 741 -172
rect 807 -138 999 -132
rect 807 -172 819 -138
rect 987 -172 999 -138
rect 807 -178 999 -172
rect 1065 -138 1257 -132
rect 1065 -172 1077 -138
rect 1245 -172 1257 -138
rect 1065 -178 1257 -172
<< properties >>
string FIXED_BBOX -1404 -257 1404 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
