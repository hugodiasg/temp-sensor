magic
tech sky130A
magscale 1 2
timestamp 1644161670
<< error_p >>
rect 1930 2716 1991 7484
rect 1930 -2384 1991 2384
rect 1930 -7484 1991 -2716
rect 2250 -7650 2311 7650
rect 2570 2599 2631 2821
rect 2570 2279 2631 2501
rect 2570 -2501 2631 -2279
rect 2570 -2821 2631 -2599
<< metal4 >>
rect -2610 7559 2609 7600
rect -2610 2641 2353 7559
rect 2589 2641 2609 7559
rect -2610 2600 2609 2641
rect -2610 2459 2609 2500
rect -2610 -2459 2353 2459
rect 2589 -2459 2609 2459
rect -2610 -2500 2609 -2459
rect -2610 -2641 2609 -2600
rect -2610 -7559 2353 -2641
rect 2589 -7559 2609 -2641
rect -2610 -7600 2609 -7559
<< via4 >>
rect 2353 2641 2589 7559
rect 2353 -2459 2589 2459
rect 2353 -7559 2589 -2641
<< mimcap2 >>
rect -2510 7460 2290 7500
rect -2510 2740 -2187 7460
rect 1967 2740 2290 7460
rect -2510 2700 2290 2740
rect -2510 2360 2290 2400
rect -2510 -2360 -2187 2360
rect 1967 -2360 2290 2360
rect -2510 -2400 2290 -2360
rect -2510 -2740 2290 -2700
rect -2510 -7460 -2187 -2740
rect 1967 -7460 2290 -2740
rect -2510 -7500 2290 -7460
<< mimcap2contact >>
rect -2187 2740 1967 7460
rect -2187 -2360 1967 2360
rect -2187 -7460 1967 -2740
<< metal5 >>
rect -270 7484 50 7650
rect 2250 7601 2570 7650
rect 2250 7559 2631 7601
rect -2211 7460 1991 7484
rect -2211 2740 -2187 7460
rect 1967 2740 1991 7460
rect -2211 2716 1991 2740
rect -270 2384 50 2716
rect 2250 2641 2353 7559
rect 2589 2641 2631 7559
rect 2250 2599 2631 2641
rect 2250 2501 2570 2599
rect 2250 2459 2631 2501
rect -2211 2360 1991 2384
rect -2211 -2360 -2187 2360
rect 1967 -2360 1991 2360
rect -2211 -2384 1991 -2360
rect -270 -2716 50 -2384
rect 2250 -2459 2353 2459
rect 2589 -2459 2631 2459
rect 2250 -2501 2631 -2459
rect 2250 -2599 2570 -2501
rect 2250 -2641 2631 -2599
rect -2211 -2740 1991 -2716
rect -2211 -7460 -2187 -2740
rect 1967 -7460 1991 -2740
rect -2211 -7484 1991 -7460
rect -270 -7650 50 -7484
rect 2250 -7559 2353 -2641
rect 2589 -7559 2631 -2641
rect 2250 -7601 2631 -7559
rect 2250 -7650 2570 -7601
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -2610 2600 2390 7600
string parameters w 24.0 l 24.0 val 1.17k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 88
string library sky130
<< end >>
