magic
tech sky130A
magscale 1 2
timestamp 1669420244
<< metal3 >>
rect -2870 2792 2869 2820
rect -2870 -2792 2785 2792
rect 2849 -2792 2869 2792
rect -2870 -2820 2869 -2792
<< via3 >>
rect 2785 -2792 2849 2792
<< mimcap >>
rect -2770 2680 2670 2720
rect -2770 -2680 -2730 2680
rect 2630 -2680 2670 2680
rect -2770 -2720 2670 -2680
<< mimcapcontact >>
rect -2730 -2680 2630 2680
<< metal4 >>
rect 2769 2792 2865 2808
rect -2731 2680 2631 2681
rect -2731 -2680 -2730 2680
rect 2630 -2680 2631 2680
rect -2731 -2681 2631 -2680
rect 2769 -2792 2785 2792
rect 2849 -2792 2865 2792
rect 2769 -2808 2865 -2792
<< properties >>
string FIXED_BBOX -2870 -2820 2770 2820
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 27.196 l 27.196 val 1.499k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
