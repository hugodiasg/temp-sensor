** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator_tb-tran.sch
**.subckt ask-modulator_tb-tran
Vdd vd GND 3.3
Vin in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 25ns 50ns)
x1 vd out in GND ask-modulator
**** begin user architecture code


*.tran 0.35n 30n
.tran 0.5n 50n
*.tran 2n 800n
*.tran 0.05n 1.3n
.control
destroy all
run
let id =-i(vdd)
let z_rlc= (out-vd)/id
let z_nmos=out/id
let z_out=z_rlc*z_nmos/(z_rlc+z_nmos)
plot z_out
plot id
plot in
plot out
*rlc
let s_rlc=(out-vd)*conj(-i(vdd))
*nmos
let s_nmos=out*conj(-i(vdd))
*ask-modulator
let s=s_nmos+s_rlc
plot s
let s_rms=sqrt(integ(s^2)/50n)
plot s_rms
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  ask-modulator.sym # of pins=4
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/ask-modulator.sch
.subckt ask-modulator  vd out in gnd
*.iopin gnd
*.ipin in
*.opin out
*.iopin vd
XM2 out in gnd gnd sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=8.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC0 vd out sky130_fd_pr__cap_mim_m3_2 W=23 L=23 MF=3 m=3
x1 vd out l0
**** begin user architecture code

*X0 out in.t0 gnd gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p
*+ ps=1.798e+07u w=0u l=0u
*X1 out.t4 out.t5 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 gnd gnd sky130_fd_pr__res_generic_l1 w=-1.40235e+12u l=2.35e+07u
*X2 out.t0 out.t1 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
*X3 out.t2 out.t3 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R1 out.n2 out 3.403
R2 out.n3 out 2.851
R3 out out.n2 1.395
R4 out.n0 out.t5 0.467
R5 out.n1 out.n0 0.465
R6 out.n3 out.t0 0.161
R7 out.n2 out.n1 0.144
R8 out.t2 out.t4 0.066
R9 out.t0 out.t2 0.066
R10 out out.n3 0.042
R11 out.n0 out.t3 0.023
R12 out.n1 out.t1 0.002
R13 in in.t0 446.69
C0 in out 0.05fF
C1 li_17191_n190# gnd 1.60fF $ **FLOATING
C2 in.t0 gnd 0.40fF
C3 out.t3 gnd 7.61fF
C4 out.t5 gnd 10.97fF
C5 out.n0 gnd 3.85fF $ **FLOATING
C6 out.t1 gnd 5.33fF
C7 out.n1 gnd 6.22fF $ **FLOATING
C8 out.n2 gnd 20.09fF $ **FLOATING
C9 out.t4 gnd 16.65fF
C10 out.t2 gnd 16.70fF
C11 out.t0 gnd 17.48fF
C12 out.n3 gnd 14.27fF $ **FLOATING
C13 out gnd 304.73fF
C14 in gnd 5.02fF

**** end user architecture code
XR1 out vd gnd sky130_fd_pr__res_high_po_5p73 L=0.56 mult=3 m=3
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym # of
*+ pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/ask_modulator/xschem/l0.sch
.subckt l0  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 1.006n m=1
Cs1 p1 net1 10.86f m=1
Cs2 p2 net2 11.96f m=1
Rs1 net1 GND 114.5 m=1
Rs2 net2 GND -66.9 m=1
R1 p2 net3 5.426 m=1
.ends

.GLOBAL GND
.end
