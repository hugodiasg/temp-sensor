* NGSPICE file created from ask-modulator.ext - technology: sky130B

.subckt sky130_fd_pr__res_xhigh_po_0p35_NVRUDW w_n202_n1098# a_n36_n932# a_n36_500#
X0 a_n36_n932# a_n36_500# w_n202_n1098# sky130_fd_pr__res_xhigh_po_0p35 l=5e+06u
C0 a_n36_n932# w_n202_n1098# 1.08fF
C1 a_n36_500# w_n202_n1098# 1.08fF
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ML7W5H a_n108_n870# a_n50_n958# w_n278_n1128#
+ a_50_n870#
X0 a_50_n870# a_n50_n958# a_n108_n870# w_n278_n1128# sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=8.7e+06u l=500000u
C0 a_50_n870# a_n108_n870# 1.16fF
C1 a_50_n870# w_n278_n1128# 0.87fF
C2 a_n108_n870# w_n278_n1128# 0.87fF
C3 a_n50_n958# w_n278_n1128# 0.52fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_EZRVX8 m4_n2510_n7390# c2_n2410_n7290# VSUBS
X0 c2_n2410_n7290# m4_n2510_n7390# sky130_fd_pr__cap_mim_m3_2 l=2.33e+07u w=2.33e+07u
X1 c2_n2410_n7290# m4_n2510_n7390# sky130_fd_pr__cap_mim_m3_2 l=2.33e+07u w=2.33e+07u
X2 c2_n2410_n7290# m4_n2510_n7390# sky130_fd_pr__cap_mim_m3_2 l=2.33e+07u w=2.33e+07u
C0 c2_n2410_n7290# m4_n2510_n7390# 108.99fF
C1 c2_n2410_n7290# VSUBS 0.24fF
C2 m4_n2510_n7390# VSUBS 27.62fF
.ends

.subckt ask-modulator in out gnd
XXR1 gnd out out sky130_fd_pr__res_xhigh_po_0p35_NVRUDW
XXM1 gnd in gnd out sky130_fd_pr__nfet_g5v0d10v5_ML7W5H
Xsky130_fd_pr__cap_mim_m3_2_EZRVX8_0 out out gnd sky130_fd_pr__cap_mim_m3_2_EZRVX8
X0 out.t2 out.t3 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
X1 out in.t0 gnd gnd sky130_fd_pr__nfet_g5v0d10v5 ad=2.523e+12p pd=1.798e+07u as=2.523e+12p ps=1.798e+07u w=0u l=0u
X2 out.t4 out.t5 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
X3 out.t0 out.t1 sky130_fd_pr__cap_mim_m3_2 l=0u w=0u
R0 out.n0 out 6.736
R1 out.t1 out.n0 5.23
R2 out out.t1 3.322
R3 out.n1 out.t3 0.472
R4 out.t1 out.n1 0.471
R5 out.n0 out.t2 0.164
R6 out.t4 out.t0 0.066
R7 out.t2 out.t4 0.066
R8 out.n1 out.t5 0.023
R9 in in.t0 448.61
C0 out in 0.05fF
C1 in.t0 gnd 0.46fF
C2 out.t0 gnd 13.53fF
C3 out.t4 gnd 13.57fF
C4 out.t2 gnd 13.79fF
C5 out.n0 gnd 44.65fF $ **FLOATING
C6 out.t5 gnd 6.18fF
C7 out.t3 gnd 8.90fF
C8 out.n1 gnd 3.13fF $ **FLOATING
C9 out.t1 gnd 58.04fF
C10 out gnd 165.23fF
C11 in gnd 5.60fF
.ends

