magic
tech sky130A
magscale 1 2
timestamp 1646019513
<< metal4 >>
rect -2664 10449 2664 10490
rect -2664 5361 2408 10449
rect 2644 5361 2664 10449
rect -2664 5320 2664 5361
rect -2664 5179 2664 5220
rect -2664 91 2408 5179
rect 2644 91 2664 5179
rect -2664 50 2664 91
rect -2664 -91 2664 -50
rect -2664 -5179 2408 -91
rect 2644 -5179 2664 -91
rect -2664 -5220 2664 -5179
rect -2664 -5361 2664 -5320
rect -2664 -10449 2408 -5361
rect 2644 -10449 2664 -5361
rect -2664 -10490 2664 -10449
<< via4 >>
rect 2408 5361 2644 10449
rect 2408 91 2644 5179
rect 2408 -5179 2644 -91
rect 2408 -10449 2644 -5361
<< mimcap2 >>
rect -2564 10350 2406 10390
rect -2564 5460 -2035 10350
rect 1877 5460 2406 10350
rect -2564 5420 2406 5460
rect -2564 5080 2406 5120
rect -2564 190 -2035 5080
rect 1877 190 2406 5080
rect -2564 150 2406 190
rect -2564 -190 2406 -150
rect -2564 -5080 -2035 -190
rect 1877 -5080 2406 -190
rect -2564 -5120 2406 -5080
rect -2564 -5460 2406 -5420
rect -2564 -10350 -2035 -5460
rect 1877 -10350 2406 -5460
rect -2564 -10390 2406 -10350
<< mimcap2contact >>
rect -2035 5460 1877 10350
rect -2035 190 1877 5080
rect -2035 -5080 1877 -190
rect -2035 -10350 1877 -5460
<< metal5 >>
rect -239 10374 81 10540
rect 2366 10449 2686 10540
rect -2059 10350 1901 10374
rect -2059 5460 -2035 10350
rect 1877 5460 1901 10350
rect -2059 5436 1901 5460
rect -239 5104 81 5436
rect 2366 5361 2408 10449
rect 2644 5361 2686 10449
rect 2366 5179 2686 5361
rect -2059 5080 1901 5104
rect -2059 190 -2035 5080
rect 1877 190 1901 5080
rect -2059 166 1901 190
rect -239 -166 81 166
rect 2366 91 2408 5179
rect 2644 91 2686 5179
rect 2366 -91 2686 91
rect -2059 -190 1901 -166
rect -2059 -5080 -2035 -190
rect 1877 -5080 1901 -190
rect -2059 -5104 1901 -5080
rect -239 -5436 81 -5104
rect 2366 -5179 2408 -91
rect 2644 -5179 2686 -91
rect 2366 -5361 2686 -5179
rect -2059 -5460 1901 -5436
rect -2059 -10350 -2035 -5460
rect 1877 -10350 1901 -5460
rect -2059 -10374 1901 -10350
rect -239 -10540 81 -10374
rect 2366 -10449 2408 -5361
rect 2644 -10449 2686 -5361
rect 2366 -10540 2686 -10449
<< properties >>
string FIXED_BBOX -2664 5320 2506 10490
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 24.85 l 24.85 val 1.253k carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 80
<< end >>
