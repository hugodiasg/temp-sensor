** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex_tb-ac.sch
**.subckt impedance-transformer-pex_tb-ac
Vin net1 GND DC 0 AC 1
Vin1 net2 GND DC 0 AC 1
R3 ns12 GND 50 m=1
R4 ns22 net2 50 m=1
xit1 ns11 ns12 GND impedance-transformer-pex
xit2 ns21 ns22 GND impedance-transformer-pex
R1 net1 net3 152 m=1
R2 GND net4 152 m=1
C1 net3 ns11 3.7p m=1
C2 net4 ns21 3.7p m=1
**** begin user architecture code



.ac lin 1MEG 1.5G 4G
.control
destroy all
set units=degrees
run

set color0=white
set color1=black

let z0=50
let zl=169

* Find two S parameters from test circuit
let s11 = v(ns11)
let s12 = v(ns12)
let s21 = v(ns21)
let s22 = v(ns22)

* Extract Y parameters
*let StoYDelS = ((1+s11)*(1+s22)-s12*s21)*z0
*let y11 = ((1+s22)*(1-s11)+s12*s21/StoYDelS
*let y12=-2*s12/StoYDelS
*let y21=-2*s21/StoYDelS
*let y22 = ((1+s11)*(1-s22)+s12+s21)/StoYDelS

* Extract Z parameters
let StoZDelS = ((1-s11)*(1-s22)-s12*s21)/z0
let z11 = ((1+s11)*(1-s22)+s12*s21)/StoZDelS
let z12 = 2*s12/StoZDelS
let z21 = 2*s21/StoZDelS
let z22=((1-s11)*(1+s22)+s12*s21)/StoZDelS

*plot z11
*plot z12
*plot z21
*plot z22 xlimit 2.4G 2.5G
*plot ph(z22) xlimit 2.4G 2.5G
*plot z22
*plot smith z22
let z_in =z11-z12*z21/(z22+z0)
let z_output=z22-(z12*z21/(z11+zl))
plot ph(z_in) ph(z_output)
plot mag(z_in) mag(z_output)
let gamma=(mag(z_output)-mag(z_in))/(mag(z_output)+mag(z_in))
plot gamma*100
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex.sym # of pins=3
** sym_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex.sym
** sch_path:
*+ /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/impedance-transformer-pex.sch
.subckt impedance-transformer-pex  in out gnd
*.iopin gnd
*.iopin in
*.iopin out
xl1 in out l1
**** begin user architecture code

** NGSPICE file created from impedance-transformer.ext - technology: sky130A

.subckt sky130_fd_pr__cap_mim_m3_2_8BMXEH c2_n2657_n10762# m4_n2757_n10862# VSUBS
X0 c2_n2657_n10762# m4_n2757_n10862# sky130_fd_pr__cap_mim_m3_2 l=2.578e+07u w=2.578e+07u
X1 c2_n2657_n10762# m4_n2757_n10862# sky130_fd_pr__cap_mim_m3_2 l=2.578e+07u w=2.578e+07u
X2 c2_n2657_n10762# m4_n2757_n10862# sky130_fd_pr__cap_mim_m3_2 l=2.578e+07u w=2.578e+07u
X3 c2_n2657_n10762# m4_n2757_n10862# sky130_fd_pr__cap_mim_m3_2 l=2.578e+07u w=2.578e+07u
C0 m4_n2757_n10862# c2_n2657_n10762# 174.60fF
C1 c2_n2657_n10762# VSUBS 0.30fF
C2 m4_n2757_n10862# VSUBS 44.26fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_U5TCJH m4_n2770_n8173# c2_n2670_n8073# VSUBS
X0 c2_n2670_n8073# m4_n2770_n8173# sky130_fd_pr__cap_mim_m3_2 l=2.591e+07u w=2.591e+07u
X1 c2_n2670_n8073# m4_n2770_n8173# sky130_fd_pr__cap_mim_m3_2 l=2.591e+07u w=2.591e+07u
X2 c2_n2670_n8073# m4_n2770_n8173# sky130_fd_pr__cap_mim_m3_2 l=2.591e+07u w=2.591e+07u
C0 m4_n2770_n8173# c2_n2670_n8073# 132.19fF
C1 c2_n2670_n8073# VSUBS 0.26fF
C2 m4_n2770_n8173# VSUBS 33.47fF
.ends

*.subckt impedance-transformer gnd out in
Xsky130_fd_pr__cap_mim_m3_2_8BMXEH_2 out gnd gnd sky130_fd_pr__cap_mim_m3_2_8BMXEH
Xsky130_fd_pr__cap_mim_m3_2_8BMXEH_3 out gnd gnd sky130_fd_pr__cap_mim_m3_2_8BMXEH
Xsky130_fd_pr__cap_mim_m3_2_U5TCJH_0 gnd in gnd sky130_fd_pr__cap_mim_m3_2_U5TCJH
Xsky130_fd_pr__cap_mim_m3_2_U5TCJH_1 gnd in gnd sky130_fd_pr__cap_mim_m3_2_U5TCJH
Xsky130_fd_pr__cap_mim_m3_2_U5TCJH_2 gnd in gnd sky130_fd_pr__cap_mim_m3_2_U5TCJH
Xsky130_fd_pr__cap_mim_m3_2_8BMXEH_0 out gnd gnd sky130_fd_pr__cap_mim_m3_2_8BMXEH
Xsky130_fd_pr__cap_mim_m3_2_8BMXEH_1 out gnd gnd sky130_fd_pr__cap_mim_m3_2_8BMXEH

R0 out out.n2 0.325
R1 out.n0 out.t7 0.1
R2 out.n1 out.n0 0.085
R3 out.n2 out.n1 0.067
R4 out.t6 out.t4 0.066
R5 out.t5 out.t6 0.066
R6 out.t7 out.t5 0.066
R7 out.t2 out.t0 0.066
R8 out.t1 out.t2 0.066
R9 out.t3 out.t1 0.066
R10 out.t14 out.t12 0.066
R11 out.t13 out.t14 0.066
R12 out.t15 out.t13 0.066
R13 out.t10 out.t8 0.066
R14 out.t9 out.t10 0.066
R15 out.t11 out.t9 0.066
R16 out.n2 out.t11 0.036
R17 out.n0 out.t3 0.018
R18 out.n1 out.t15 0.018
R19 in in.n1 0.704
R20 in.n0 in.t6 0.124
R21 in.n1 in.n0 0.096
R22 in.t7 in.t8 0.066
R23 in.t6 in.t7 0.066
R24 in.t4 in.t5 0.066
R25 in.t3 in.t4 0.066
R26 in.t1 in.t2 0.066
R27 in.t0 in.t1 0.066
R28 in.n0 in.t3 0.026
R29 in.n1 in.t0 0.026
C0 in.t2 gnd 40.33fF
C1 in.t1 gnd 40.42fF
C2 in.t0 gnd 37.40fF
C3 in.t5 gnd 40.33fF
C4 in.t4 gnd 40.42fF
C5 in.t3 gnd 37.40fF
C6 in.t8 gnd 40.33fF
C7 in.t7 gnd 40.42fF
C8 in.t6 gnd 36.14fF
C9 in.n0 gnd 10.99fF $ **FLOATING
C10 in.n1 gnd 56.69fF $ **FLOATING
C11 out.t12 gnd 39.58fF
C12 out.t14 gnd 39.67fF
C13 out.t13 gnd 39.67fF
C14 out.t15 gnd 35.25fF
C15 out.t0 gnd 39.58fF
C16 out.t2 gnd 39.67fF
C17 out.t1 gnd 39.67fF
C18 out.t3 gnd 35.25fF
C19 out.t4 gnd 39.58fF
C20 out.t6 gnd 39.67fF
C21 out.t5 gnd 39.67fF
C22 out.t7 gnd 76.39fF
C23 out.n0 gnd 22.95fF $ **FLOATING
C24 out.n1 gnd 13.15fF $ **FLOATING
C25 out.t8 gnd 39.58fF
C26 out.t10 gnd 39.67fF
C27 out.t9 gnd 39.67fF
C28 out.t11 gnd 38.21fF
C29 out.n2 gnd 42.74fF $ **FLOATING
C30 out gnd 59.84fF
C31 in gnd 44.14fF
*.ends



**** end user architecture code
.ends


* expanding   symbol:  /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sym
*+ # of pins=2
** sym_path: /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sym
** sch_path: /home/hugodg/projects_sky130/temp_sensor/impedance-transformer/xschem/l1.sch
.subckt l1  p1 p2
*.iopin p2
*.iopin p1
L0 p1 net3 529.2p m=1
Cs1 p1 net1 29.38f m=1
Cs2 p2 net2 25f m=1
Rs1 net1 GND 69.31 m=1
Rs2 net2 GND 3.196 m=1
R1 p2 net3 2.702 m=1
.ends

.GLOBAL GND
.end
